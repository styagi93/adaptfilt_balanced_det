��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[P3-L5���4K\��q��M�U�}A4�Z�MT�����~��h	)��6�!XK=��HNk$���"���O�-�� �_��a�g�/�[�6�� KRӎMz{|ˏ���'�3�2(�.<���( ��I�F��^IG�|b�d(��1�b�D�^���q�17a��1R�u*3�������{Jmy������,����rn�c��0� �0G�y1�i�8؈o3wO�qvY�Ե1��3����kD�#G��~�P�܊$&cݬV|"a�ч�n����;�L"?�J�7of��_?%������g��Y��
j�쫈��Td�0��P�F�q!.����z���¡�j���w����DZ`{�@Hxn���x	����2,����|5
mc%N��ԧ��5�5�?r�k�T_��ƌ���(�[$�ފ��a��.�E2݉�4$����}l�w�x�q4B���l��b� k�(�e��l���Vĳ�D�ܽ�n���1n�)�LV��Kɒ�5涰������DEɣ�, ��L9��_�R�J�3��GXF�j��7�����)�Lx���U�������:=%�`�7�T�K�*�7�K<l]���*ƎfsgX�}��a8�G��+=�˾�,��;I�O?ࣱ��zb=�ku�Z���%
j��ڂ�s�����ϫ�F�������-�$m�S�jO��b�]����}M8z�V�;w7>�<R�N����.�)�g}��� �?��X�H�����c�]�]���1�(K�\=\�7^�	%�l?�p�� �L� AIp��hA��c=Ie�JhE����#nF�Ӌ�ϸ��(��P��<�5&�B{���KKll ��y�>��L���{�*�)S��+�=�k�V�k�ڪ� �P����^�̊��a���*�ȿO��|�ޏ(4��"��X+��Tc.�@��T`=�jy�i�a� ��PpU���;��%��n�vW( ��<!���� ����H��1셄(�'K/�3����*[�k�w�h��~��`��Jdٞ����Kj\?A�k��w�D_�)�듬�G��&l��,�M�j(P����K�g���=���#�'�v���K��;Au���qI��A��+����~��E��ϱG�{�t�G��1�d4K�Q���F={�)p�U�|V��%Nq(�ƈ!�I������!�n�"��֋[M�)�y��$8Z9��A������ލ/C�iY�o�����D����߫�е�{�H��g�գ۹�d�u8����eeӈrQ����^���w�G/8�O����&�0�F`Z��'bs�ڜ��ޖ���`�R��FB�C_��ّV͵�H����A}D�V�)	��	�V�����1
}�Q(A�}���8�a���t��ql5ɻ`=��iA�8��j�CV�3@�=+¬�L�x����̐E׉��Ԉ�Z�9[���1����t�نgj��+�e��oR�ۊXE(���.U�`�Tp��u��=���^�GxUzz�]m����Oktb�BT�،�t� Qw��7G�1�?v��x.3UE�"��Y��}��n!E1 L�RKI�@��\����O���P����2u��iX����;�U�F���H��m�:�vq��das�&����k�
�����w�$�`c7��{Ek�����F�o_��_ɴO��u�L�g}����I��ZHx����83�󝶿��,B(��db%m��EFČ��&=��>���DVc�´byV�bW#!Qքܬ�$i]3}���>qґtp�O�zK��F����s���Q������l���!9�!󋂱s��0�jWp���I��'�[�#�`4ܬ��ͺ�H� ��A(k,�8�"�s0��^������$�(�(��ľ�E0Ŋ�|��u� �臼&<�J
�D� .�;�)�
�ۧ���ʠ6�췑�v��K��1�`��!�
����x_l�AY*2]�o��ls���ˠ����N�����:=ƶOVrt���3�f+��]-r�}q��d��l%Rs�?�ʇZ����j�%��{,]�{��W��T���+y�|U�:L5Х#K<Խd/T{� �ܠ�����1�pBm4�oi�o��K�f6�s{���]>س���� ���?V��3��x�n͇=|�>�mɀ��K}�6f�7&W%�/�Z�ǑN��U��'�a�Ҿ_���h�W6�a���bwX�w�,�$�@��ۂ���r��^
�-��]���'Y{=0L��~��l FHr�DV��')��͸��g��dAC?��:���3oN�tt�Z���B��>]F�a�"y+N��͍�ΐ����$4�J�^N�UXJ�����m�B��m*��6xP��|yʓ@�6��4�.����Z��׼�dڝBìUg$~)��	,�h�="п>٫�dw�K�S�������wk�}�Ĳ�������LPVr*�C����8#�!�E)�k�4++26m}O�зzSeM���l<��%��?jCUVH�E���h*!�AP�q���)UD�0j��-I[Z��zB�L�O�P��y��6x/�	K?�2���k�5���8"{�|a{�NT��o��]؎2�a������=���f����'�z�9�smiJZ&E$�o/@<
9�F�.MA[�#�=ͩ�σP��b�04z�|����pK�Djl���ixғp��H5�^w�D�Z<�@.���/�����oꃪ"�����W��Y�0�����WTv��ͫ�K5��a���;r����	�RT�$n���Y�ý��\��#����������B�t����(�����⸰�E���Ҡ�FA���u��ӪN��P�=�X�~�S����:*'�0�F%9۩"Y���o"`Y"��ֹaW&Y[�$�����{A�TAO��݀�E�N}m�^����ŗr��$$�@���[%[���F�r�ڮ��L^%�
����`IH����3���3GfS��r���������c,35Џ�fh[Q�%��os�9k��'��G�M>w�jV��a��K�?����ۄ�8�ԇQ��E�����+�^�._���|{��5��qu=y�Lp8B\�w3�����Y��6W�	~S�O!"�H���SL�Uݤļ+D��MtF��WU��yZT��ѥԮ�D��%IZ�ڀQ$9T!�8]��{CY}���}epHN�&�	4��%I�W���B�r�)ޫ�Dt��P��ߵ[�����L��^�f`Nl�*���<%Y�:�U	�����%�Ld妀��hg���*��
�W������m�a�� ��o4:�"�9�Y�|/�B����˷M��!㨵+D�������%�i���L��W��>	B�\ĽHv�)���-��\��TwS������8�z��D�_��c8�v����I�������x_����x���v����)�	�/h�hl	vg]��$D�����{D��<W�Ii�T�z�����ќ�0Һt}3�b��;?<��-�ļ$m4q/=�#����~Z�B�7�s^Eu��3(J��b��\#���2_��L���>%�|@~P23M��PTX��|�Ή)����r ����R���CYz�!��<�,_Z_�3�G��w2��Պ`� �3G��uM��#�Z�>z�Rr׫ď�F�,Qx��Y:I�~,�v��QXH��gV���_y�h�.tz���Y�"����޶c;��frt��n5
�\�0w,lj	|��W�N9�2�>g�eR����d����<�k&�)ɝ�M"�bk���CBߴ|T "��Qb�;�ZV��U�������ZI'5q��+J�檀�Y��\i,���Ќ](�e��*�F�2&��4����1*Z�e�:�Y8N��R@���*�a�B}�'�D\ѣEhy��,�=��0q(��b�]n��t�������T�0�	Bw�i�ynU�����*�+��Uj�d���Ȑ���C��.t��4���{N�ʹf������շ��]������.��@�������<�D�M�j@�w�urs��9��>᳐��cO�ܲ�O��kɼ;�*!L�����jl�_��b�B���pɅ��H�*jo���elfc�e�ha`�R�+��.���;�L.X���a�4���ד��x�;�B>��j*�j~ٲ���fY�98U(8�ɾ���N����E�����v:�4y�f�җ́�+���n ;
�&(8i4��ф�~	K�'�D$��j�a��xQe;��s�+����[�G/\Y���v_U��x�Q�d���+�{х���1�H�<iX�sLW_���"�O�� ��!��nW�8�U
��˟��LE�Z����X�m�i���J^Ds�eh�j�72R��=|J�I�4��i�Ln#e��,?�oagɀ3b�0�A�H?��}V}�ڢ��KO�'�W��*�H4�
�N�%���]�B�,7�xX6��{��f����	�"��U �ؐ]�*�K�����@�TL.G�' ��N]�z2rV4)<��9�iv�!�DI=Ft<2t���&Rx�Z�H�D�pE������M���g�A�J�;�|!�H���(�Qx�lfKʁ|�q�����C��Ѹ�����!C�Fo6I�)��q<�̄��.U�w;Z�]eu�����Z������{�ڐ�(2T�����!!�6Qu��m�%&M|l3,�Ă�jf1t��2��s$_.��q1�"�(��{�G� iB=HeM�Uh�ז��!:�P[�S����H�\+�;F���U#��sڂ�+E��h�(K?�ps�wа��t�L ����o��'���Étٶcg@Rr1|3�z&>��^Y��ϫ�t�7#W��5V*ʼ�z��M/���1��{k)=mD6n�T�o=�C�5��Gn���1�F�eMykι�cg�at6 z<[��ᆜ����1	V�Δ�
��,�j�c&����J�����Q,�I!-���������p�rv�	ͬ��� ԗ�.�g�V1��D���t�p�^��P(M�'�;����*�HC���NQ�M�:��D������ܙ�a�k�����A����rx�J��^qS�e�J�N|��\�%��wnA�%�,���t`��o0�ڒ�QY�E]��a5�E�*֢�Q; ����d9v���c���^����	��z�|��ݵ��^�ȱ����4}�O�1�.��3ʘ��P?j�a�X�9�	秾�p��"�[Ol}�L��`��=[Ս'L�,Ɩ�a��7�hv�rv�*q�MP.1�����	)���>�j�;l5��@p��pGp���j'u9M$߂TlD$��1ԈA�hy��$�%��;�]�[�.N���^��.D���X�UšL ��~GN*�����YXR��p����s�ξ;j�����r�X�t|m��.�RHj�ɵ#+�W�� �*�g�yPm�U�x���3��<��P+uo�p�-9����I����,�
0>�48�'$z�I��`j�u׹�n�mz�09 l�X)��<��1ˇ�$j���BM����sJ��/2�Ρ)�ś�Fu�iB\�;*�Zy�RfڼA��c��N�Ft(��v�e�������HL&	j�Tk�����}?#A@���~棊��K|E�Ժ�e3X�lCF��^�����l�vT��}k��R���l	`/��:�<iʫ�2�>yS9���e�����݋c�ZQqpĺVΎ�u*˕�W1!�1f�s����wb����8[q�fN����U�*�Mf3Ie�����������:_hに�S��Om�U��e�>\�kҼ�i�/`ӫG�wM��KX*;�Z���s\�ڨ�OlR�`@�tߎ���c?t��!ᕂ�f�(/]kL̚������'kDm�����w�9��5[��m��G�E��0�ҹr�%P%:er���j'����%��d���ȓ-��nP��IGמ�����Fy¾iB8�s*�s
z%���읣�=�P�����)|���@c� 7\���"��5?C!(SP�Xy��9����}��r���� �*:f"�����"#d���&e�C�j���-ף����b"g��q�܉�B$z�d����}:�(cBIh���T2���.���k������ 8d��-��ߌ�f-&�G���J��!u�H^+�z �E�1˭�����D\�r	%����0�(��V2	k�� ��?iI7�R�NEy	Qd��y��q4g����_D0_x���7���V��u�a�hx�5����몂Y�����-�^�p>Cڼ�d��)��<ܠ۸�1R�:<��J���*N.�2�)���p,�q�sM�;�T��ݕ��.�f_Z���r2 ɲ�S6@�Y��DG��� �6F���������u��~1*7��� Ly;��Ĭ����*tWʹ.�K�Xc��X�fO�a����$D�\=�8��W�q�^��+�+��E�R�z�z^1��@5�zQ����:�c��Y�P��_`�(��\_�d�戰A�Φ�s�&Lz0��E������!)�6�6�|I���/�ʊ�3>�t	.@�qʳ6[�&���'�~����OR���x�*���fУq��te�j���j������;�?a�H��R�Fnm���g�yじ��5C����\�pv�0͝_�հ��,@,)�����[R���� ��;��?.d_�@�[��	�g�'���{��HZ�����ާ�aLOy^;�1�ڻ�gA��p���Lˆ��H@'t |�hZ��%���#��&�L�U>|N�����5{�W�[�Q�Q�Y_�%>����&}yiƋ�o��9A}������bf~B�� ��K�&(�Y�I��IV�t��{_�Ç�~��2R����ҀC^�IlA�m�o_�ʀ���j��Iy2��S\<�A��A�VCa6A��Nx,�ϓ�$��܉��00�9.�L�ZF�I[R�ؕ!�^8��Y6C���?�iOZ�,�,�{R>���7h��d�`۞L�~Y 8?�v����3�~Mq��u���3�h��K-ș����G��Iέ2EA�V��FOjh��1��lC�_u&���.��%��q����"�:���lI�˖�������<�w�zH,���Ｖ�!m��}'c)e�]���>��yǦ��R=��@JGKG�z�ZU�6��0��SOD�_kp-}t �|(��g��;�I�ֽ�	����t�jYo] S���J��w��R���4[�nH(|(�ڞ�=�r�ٕ��x$SH�[O�B��0��̬�0ݕ�#x�
��3�-KH�%	x ���ޥ��\9������gc�����C��E_	�����(�f���"��u�m���i� �������B�,�H�����ƽ �s�%�g%�M�R�p���CO���k���'��H�;��{�Z�xH�17'��_����C& �I%`D&$yu�x*l�e���A���j\����H��l�^�E��Cd0T��ι�%�b'��Ĝ)�YX��Ⱦg�a�A�FM�94����#�k�9ħ�W��pM���U@��|���XD�^&�P�N��a��P��Ӭou�X��N�}��C2�]���o�7���]/
���P��#��tU�bl�>��X���b%�����C�5⡛��ߜ�-},��e��U�1�Co#�WJ��UbHC����"�O]�u���Ø���jg[	��kX���2���u��{rt��K��c�ޖ���ă�w������ج�ޖ�X���<7|8z���d秊���߰b`o��۳A}+x�W�u��H������%���[����)o����=�{{8�_a2hAA���eN�L6PA}J��[/�D�/�z����|�a8e�"��6>��F��a���q1m���%N�V�@�U���W ���k�6�U����k���Wr�-���F)'�b�F�΢��2�pb�'2w-r��`!�亜;�8��K^n���o�E�׀�@��W���剈�Ucj���NTl�rFL��0K��a��?=u*9�*�A؆������[8�L}Pw�l�/���Ë���?�� ���T&��v���u�³�O$ޡ�P���QHW��n���y��߲QE0�a�|�'�:��hӢ쬧&r���h ����a��G]�;G�pk�-O����8���1�`��C�^�S�o&\�\���ly�+MǉlH#F<U���j�v�'m��U�3��x��O�bu�ԥ���K �tYV�r�e�&�ƹa�r\�Bȩ��á���]��k��+O�%�}�m��@������Q�=��SsQ�8G�z��m�ye(����@
^�7��lѵ^2�Ǹ�K���l�(v�?�ؔS�=p��!Q��R�Db�&$~���/���Y�[J4���&qХ��Ic�/rj�(���:&� ���TwY 4��"#ns�p}���q�� tԎQ;U��J�R5V[�h���֠���5TkqG[B���Ģ!*���Y�ڼ��I��W_n/���mx�ӖIMq8�c�!n�\�(��\XS��:�v�L�B�`��t	 F�x�2�������0�'���' 7W���>N|�~a����,���$��} '<5R�
'���֍�����,x��<����� ���U<K6qov7{9�^����[��-c�d�����-�թ(�\���B����zշ6��D�z,?sƹoM�nM�k:��l0[H=\ۻpIp�L�V��{
��a���4�@�1�}-p�f�T[Ei!�N��tR�w(ycO�1������$S����z��:�@p�(�<���Պ�Q��ƙ�jV+���d 9'���@nK�R/O��,/�Q�&x�7%�U���:�ؚ�3@v`QnC��l���4R��i���|�����R����k��_�¡��-��p�q���!1���Ħ2���Q�?�s9�!"F��=E�K�>���&��w�A:���Wl�2����1_t�p"���za���v�֓x5�t`-fVVk{>��S��r�/Dn��p�rm|�����Z�^x��褈��h*�!��C��Ƞ�c��w@�`bu�m#�#��T���
���¤ܢ�-��W,�(��E8�$��j7%u�;ۆ]Q��j��\dƎ�b)�_�p�#�4���7W��l*���tz��Su����t�xV\jw�����V��	�i�Xye�w�L��2�q���A�t�k�X(��͖!ȵ�"un�%���v[�v�+����b-����l���0i�ih����v���q��?b�����'�ˣ^>�)���`�l݁w�-8�`�	�"\a����-˺�u�������.��d�E��Zp�ހ�T@	&�Kai��\�F� �B����;���_�,_@�3��(|��6���O~ap�%W�%��r�3������k��>(�	?z���	aCfx ��)��;�I!x����$+5�e�W��J!��+,�6��� ?Y�f���t\/O�>Wٺ#F�L�BtH'�� x&g
(p:t:N�P���Cr����]q�m�r!�'z��d��ޕ�(�o=�}�ض���O��DV��MOy���tǁw��g,�ZͰS�����J&5[��n
	�N��X�m����^CR�Z�=qD��ĳT���������Z�Ì��G�yWC���$�2�_�c��ŧT�n����dE��(
Mp���%��g���EC�$�^�X��8G�8���+��$EΣ�-�Sid�k�Ʒ����c#�Yi���+�RL�n��euBp/�c?�zx���H$��*���iG����g*���Dn��~�7^�
�t��erkX��˨�p~��G[F���?�q5e�ozk�;E?�n�?�@������ �L۞����l��P=�͉#�����D�Z�� �J��+W^����c��.��JRz�v)��m�e�J�XQ�X��p�G6ێ�c��C'�k���?I������0/e�;�m�5�W�}��73ue�*+��/��p")u��#8�	�IR):XrE|����/��#���+�%@vt^�{��4F��T�}`ȡn��L��f���o@Jq�4f�̝�x��@�Y����1З;�1_����z)��!b����J�NZ ��="�Q҃�Τ&}*���ji�?�8���41*��	��gן���S�|ẉ���潆:���[�����Y���e_����������"A���70ܪGB)���i���8* ��c�A�]��<�a�b�y�<{w�P����y��w�!|Cg���Ո���d�q�e2]����-��ߛt��dґ�	�|v��X6��n]�^^��{�[#�45/5�4�Nʾk= T�ӵo&l�i��R������6cd�#�uc\�;@�NaN�a\I�C��e�~B��6��],��=�ꗱL�e���Tbm�m�`/��E�Eۀ�
���$|$����g�cy� � e��Gv+^�D};/=��x��9���W��˫���iUQ����g�C�8�%Ȳ�:T�ś�3��7� <�/=��s-Bg���dV���H�k�wt�I��K�Z��������&�c��>�nR��x�(����aAF��J"uȒ��J`+`�(
�������'��##����u0��QB�Ǩ+��H���hҩ�էSs������\�����x�[#��*\!��f�?+l��1?�)���Vʤ9�������j�3���#�W�2_�焔����I5G��A�gԺ���b<��;����	��WB��+_�@iH\��d�<���#M��T"�O�o��&K��*���D񁺳�1=�WC9����Qz+M|�9��96�4k�I�U��h���%�+�ς�5��xw+���<q*�p��t��)Ȝ���X�n$��E&y�*>�G-�j�?��.@�ex��Nhˇ$�%�/�4�FJ�W�#:��57IEL۵J����UA��Ǝ?V{]-�>��r���}�̶�3ϛ��f��7�s��!�1�EÆ�:XU^)|7� a6�Ja�N"Z�K*#WK���ϔ$��[z�y\p��6��	8b
s����mU������r �����P�M�1@N�y�窉�,���MF�CF��E�Mյs�|�9[́�3ؕ]f�]/��$o�
8yp�44G���a�3(��6%�KW˸���^�e���	���V��]� �����z��l��'C�(nIh�t5�釃9���
���%�͔��i�l4��t�p6.���4�{���p��vm� H��r���FJ�i疗nʴ�ѣB�ı�Fb�O��tV�U���Wf�[��ġ��hYB�\��8�®JfaTd*���#�1d>�1�'b�9dYѥ�*V��6����y��o����i�����s��u}A�e�P�d
��SY�����U�l'.8'�&��N�m�2C�w۲��]���+d��	O?��d|�2���Z�ŵ}�6u���/���N����ޜ� ̌|�(�f��"��p�ѫ�N{�W�O��q�'��I�{�����7�O1�%�zI��t��YHǭ�,�I���(���A#�k���r�l�r&�wH8�G�Ǽ�=�F�)�4�?H��n���ʝ�
˃�N����
�}��k2�3xa��P�C�`V@7E��d���k���#k�u|��5m�}(c|���<�
��v*ǘ�S`��Co'v]#�h�V�&��,u<,����>0;�1��%1aR�{�,�T�+]�d#�/C��U�n��e|���HK(��˼E���g�j�M�����xK�jb��	����tj �8�Iw@`��3G���W-�2�k�����l��� ����Sח��7x�?�W����/8K�ڸ�Q|g�����S��\^�S��cvC�⍱�aӲ{w-��Z*[�Au�Qܚ��f&����n��NG ��Z��O�0�Ev��B�W�O	S��K����"a3}�Ϙ��Nf�/z��z��x�
?k)4MfL���K������E��<<b��0������S�7�������O�k�殝���jL�`"��9�ZKp8hM�t[{y�|B(VbE�˶`��B(���ۏ���1G�k�Ը��7��v܂�8 �>*�1�|j/�q�ށ��"��"-�s��kd�s��?��B��)�ʂ����P^H%��0Ds��h�M�d,�0t�I�4�<�h�Ä�{`�ሯ�Yfb�.�Y��6�K����x����bu���*@���
ݟj0���RK��{���������;�V��&u)�'�qO��6�ba;�s���[q�vW���yD��b�΢�R�	��Ik)���7f�+����e1)�T����$���$�=%����.L�)���������(�>�2���L�+:S��x�c����ٌ��Z��˲;��d�͔�[б0�ƍԟ��g[�8k+[z��n��E�߿����8���lf�|�VNQ�1 ��PvՄ\�i��i>o]r�`+TF�	��Ʌ�W�i)W��a��D��־if�(M_���E˱��O�t��3��>�&)���t�rxX.�6F�s���� t�d6��\�����z`(3RP�`��\��~�z�@�cWh�ܖu��)�����9W�wE�C��i݊��/�W���l����u�ٲ��������dM�m�Y�?�n��Q�N"�O���N<&�i�G�*���sc�s��ې6�����b%�)5~_���u3"�6�W;(.QtH<����+���0�$lC�����-���T��H��q�{\�RU�SxD��xr1��"��pۥV!O�ʗ�|�ji�B���$�ߧ[m
��p������H/&����x���&��𳶑,���W�a�A�g
o<fU�5�AR\��8G��b!M�- ��aG���.=�њ���[C��I��o�t�=Ryߐ�EL����ު����V=un�ug�u�%Q��/ޢ�~�I�$T�wP?�RB�"o+5�r���B���8eYŇ[\��d�:��zX'ҞA�1ƍ�"���u�-+G-Q
c�"�Q�����o�!���j���aϏ��f�j� �ԅ3�$�R3t��ֿkv��5!b}��1>���^�5��:0���/�~au�Y�1��jb̌�4{&�E�\�
�L���懪�"�7I�	*Bڦ�	���n��W�~L�Z��_)U�4�i�$��4q�w.I����r/���ѧfL@U�>9@�E��3�T�*k+f�-zS_h��36� ����jZ;��ρF�b���hU�*���N=���K���T�ͬ;]+FS�mP����m�&5P��xkq(�Eѧ�����۔T��-���!�iJ��4Z��VM������1�Hj�,S�	�w�[@�X[l���C?���G�Q(E����]N��z�H�D���!Bɽ6j�^ГC<�m\C$o���f>�x,T.�]/�Uo�}~=�18+N��bڞ̓E+�{����w�V�;�'�R��)2;j��
X�_����3g�5)�O�Xu�ҧgK<��@��̊�-����@ƾ]x�ܭ��?v�4��k{T�1��T�7�X̑��:��b�i����\�3Fu֊Y��������B$��
>	t�L���`�v�l�ޙ	H��42��.�g1�3f�m�!
�
,�N��$g	�.D��0��N�}O>�fƥ?�\�Nn=$���T�*�i�n�'"Qk0�GoC�W>�:����.�L�^�.�E�g��wY(z<����ee�z�|s�u���}d;�I�W��G{@���=��ڣ�?HS�����Y�x�
��B�O�a��]�G�/�\d�VKy�{����m:��F[�jI�4�HC?-����I�N�j7^�I�A�.�L����-���2Om�K���uD�2<�R,�U�Hη۫�� ��q�l
��M==P����߬�.n	7�N5~Q����n�۷/&��x0m�7TR�!����`�_�WN��YIt�3�q������z��l|�CU*sqhљ�T)l�XM�ӿ@W�0�j)�w詙wW|� ��|���a�H�bN���||�|ޥ�f��x�IԶ�����{��(=����8]&�ݦ�A�(�x���/�;I��y��P=�n�8��.� �h�cZ��l��"�I�>�5�?Υ���xh-a7���QG���4�VW���"�xcs��G�٪�m���,�CK[�0!6�j��7��q
t¼P��W�i��F��PJ^T��c�O�����t����9M��T
���xP�滖at�E�mWX�Sc[���؋~���k�l�O��8 ��@�^6�M�p�å��̍�����e�q<�b��QOMʶ\Ch�����3Gu�%��#�@�Ė��"��
�)�"�2�TT���8'�-6�eC�`�&�P+����)���uyغ�թ(OPwvnப,3���ھV��`ԝ�qN�y��YϹ��Z�q��h7��4w�x-���K�`Pj���]��3�d>+X���-g��X�P��.H�1W$� �WzR.%]��W��O���֏uJ��e� ���g���v�:�`����`�d��/gt,[
��F�SI6� ��~�V�dÇ�_��F"墚�Ec��v��>˾�)�-�ѷ��T��-)g��;�CZNY��il)ښ����������F����s�.ф�S�j��[N.���6���/��*6*�.��H�1"�N�B=	\܄S�K��ͅqL�f�ȧ4������ .,I.�~I01�B�mo�Y�u�b�M�v#����ӯ&$0�8�X�lN-����#��J x4�F�#vL^��r[b���DBP�v���A��*C�:��᜼���"��Eӓð��(v�,͖۟��Zk&L�of5��8�d����+J���\�ک\M���؜��C;۝�iT�ͣ5�v��q�}��8��~`�����fb��XCWw��|��h�3�����*D�@�gJ�w�E�����^J҉2%�$���4�4NE�ڐ��Ѹ��6�Gp+����2�$q��G&[O��B��ɉʯ��LM���1O����ga0��^��vf�Е�5b<�v������ҹvi�'er�y�;�۷��KU�h�&ѢT̑2��[h����z�I�/�{�]o[P �p���\�qb�1���l�<r�V�O��p�/���\ &�I�!��(H���FH���t��4�N0���{@�K�6n���C��߱�P�;��i�F��r*�j�*-Ӂ��+D�G�$����k�+I���6��L��]��\�a����<A��Y�=���Q��m����\^C�+��i���+��B�-���A�-&=�͢���}��ݑVx���I���B C���6%
�C�����ظ��W������U\r|/!_~$�_�|b�55H�� U<r�I)�t�!�$;�A���G
o�{����3����(���΄|-)!~lgM;�t�:�?xTO����|_��az\��?��:k�C͓͵>��73s�6@Zq�q���k��3g�Ƒ�����|�sŹ���C��������8����bRyCS��Da����|D�#&�9�o�Y�OY�::y���{t |��H[��T��V�d�(�饄@��3�>�Y�˝�C�0ь�nI1�,��Y��o�Z��������
q��ۏeLm't����g�Z���%3踴�	�JՎ�Y��l���E�KB����*���yKđ]5���K#�b��,�O��sf���B��_B��3%/�A,����$(��/������0skf���}�B �m @��O�>ƶ���j�ܔ��[ğ�r�kB����?_37��z�[�m� �Α2aT�qͯ�mG��t}���hkU�%5kilr7\[�R1����ֽ�堑�	���M�ڍҷ��b��S�|����.t���%�W��������x�\>>2T���=�=�O�����s'��=����122�������CE4�����Dsv����.���{�ȴ�
&��,#�[,��7��}��?�1 �8�.�2�)���vD�9֞/�@���	eSΩ���Q�]�27}OϲFR�w4�H@��/t��n�}��|�<��v��I��㓲&�9�G���.�z����q<EZݟ�'ZI��ۏ*��J1�{°~w��]�X^c�~n
� ��J
Xs����m5�#�k{�^�E�H�!�N0�TCU����syE���5����̐�e��� yx��leH��gҴ�r߾$&�<�
atA�\�/yė?��Ӯ����K�9ˡ�k�G���p��6�����x�j�AxoAt��h[m ���P7�;.h�����u��K�ɱD%��ʂ���P����bx���>����RC��E��C���1�0K�ڶ[l��:�<3��ى�㣢�Q���/�:�kP/�{�	� ���W�U!ئ#��/�T�|��qdO��Tqg��`��19�tU�G����,�~�ΐ�w��>�㼭��C	E������/���,:�'ܥ�x�U�j�^����o-<$0�Ȑ,�\�j�%�>/��uhN*VX��+՚ٔPY�������_5�E���~U��ܨ�]N>=9�Fz�>�d��!Q ������5�,��0W5�Vb,�Ք?^PH�[�&���ᘙ&|�5\1[�;��J�3y�����l�l�b'�'��EΚ!����
�zK�pڵm�欮LX*N��u�d^8���f��Ow O�D���)�T�D������l�� �4����G4�3: P!ݜ7�DP�fv������h��G�߇;��^Z�qp�൙2��(��vJ�a2u����C��RC�A%���Vg,�'��U0H@)".L�����f�xk�o���lOBP�B�8�7r�a�d ��EB�+Xf��n�_J�����J�VoW�����#��a��Z�L��Uê���XP_����WG4% ����K�1X��o~s�K�f�K���Y��Bd$#�v��0p�F�,jm�S���'��[�g����1��N��1ux���x����)�h��"�
�l"=ۖi)B`*?T�D���M�
g��RY'?���A�^��I��<�rC������ �V;0�����wK��4g߻�	^�ӂ��g2X����,�EZ1ᆢ�������`(�B%��8�?��71p
cFdD��4����l���-�3D:;f����R�;G�	��1E�P���G{�K��]��&~�s�R8�b}�*�0��X��//�qi��e�;��V7��ƧF�s,0�j	����p�VHC���� v��o4�������1�wU���v���*�%�i��!��n�������d��A��_�Ml�sS`��7,�w	��s�ߑќ���<4E��2�H)��Y�[�<��R�u�mex��?_�
�7Dqy?n��`%�O����,Z0��-���B��d��$�\7g��`B��(:zv2���5L��:gO�]�v!Y�
c���[��Ï��; �yQp))z��9�m�Yķ�w��{�ɞ�Ց�?���V�[��� �2(�j��.���O�&���{��|�rn+%		߁�c���O �Kj /F�m��Z.�5�C������
��/�K�@B��i�2�<����&ګ��%�'�A;��Q��W�'�{�G�2G3[d����9�B�0���ިdZs\�I��S��J�4�`܁�t&��}LW� ��_�޽̘������Bwea�5�;N�涧vqѹ�>����]��{���; oi�K�*��_��>Z, ����#~s�H�l����S�
�kP���rr�xg�!�a� �٤��WҐ-��&�91� ��[�R�\�����,�U��I��+L���/=�b_ckJMv}R��6Gܨ;E���)\�DGءv�D�{��NJ�f��\D*�:ix]�Co��[�QlPZ�y�#s�Y��o_Qc�$ZhVk\�p����ȇ�++�Zn���y��6g������+L���e#���t��`�ȿ*�'��l�k�j��H�s�bZ?��X���:J�!���ȣ_��w(8������o��b\�V6�������'o��ZiCq���36�R|"���C���R�@�/v����VY0�@��"���G'kP+�:�G�������J��mr$���4�[�l��rjy�nR1�#��>��FM��,�²V���m-�gʵ�\?�+�0i�޳4��2�P&�E��f'��:� d�VĚ�$BZ�G��"G�N�6�=pNq/Q3����VhT�ɤ=C�Rӣ"c��ϭ$�X��yU�����6)�g�}8*2�p[�#"�8�l%�(��p������#���y�Y2Cz�b�|��(�4����B���O	#qV+~�
D>��7
p�n�z|䣬`�-q��qf���g/�<�����XN�y,���]�F�����~9?,�N�?��.21���܀�oW���� 4=}���$�53��a{˻W��ϩ�u�Y�룬��k��`�fqd�ġu�gO@t�#N�	�#p�9 ���S��j��`o�#��j[$�K]1�����^���x�J����J�r�b��RNC,�����-0W���*ܵT�oI��`�Ұ��,y�5ax����:0�-9H�8	���f�Ք�+$Q^=�?P��.A�H��.q�>��<a��0����)=��|���������o�N�p&c+�|]���<z�����#�e�,�^�1�%#kq��̖H�	����l1QƇ���ɇP�j��|����̝2���y�O�g��q��3��������NY����11�2m�r���4����ca\�T�x$ >����"q��4K�Or�95�]V���b����v�!�x���B�QgW����mQ�T�It�
 �"�~��rm���7� ���#"|k�2�|b08���6"No�J�;�J`-�B8�6D�Jsx9����V#V�=44���t�m΁�sӜ����+�F2��k�k}G�aaّ~/�TQ�5‧gV�X(�^�Q� �4��k&����vM8����4O�G@s���X=� q����7���:�Z��u����6+(��K�j�ZQ�#�,�9��A��S��5:]r�X��-��)@�Q$�Vl��sl�󽼝^�=��N���G)j�LE���Q�<��	�lӌ�C}�Ӵ¤������Ӿ��
,��k����A��΄2�;^ ��������ǩq�;���/���~�����"���.�v�jA�֠�,����d�l����������$����=.��Gc�����o6��-yR��kܿ4�v�Q�E�we�� �iԸB� ��c�C]��Fk�&4M �.� ���������Fˉ�fyI C�|p��yn�[�quQCDÕ�}�`6�T�I'�y�YAN�x�"�dF���(����4r�0��љ�_㻮�gb�u>텆�~(���^�3M '�p��/��+�]�{�� T�a 5�/�=�n촛,b������\C�yX�O�'�o�s��'���.� ���fT�`�_-�����E�W��4Hr�]�cד�0+_��t����f�Dd�IY����N�}R���oTKC"����(bK� `p�-��1����y	%*����pnOd�̽kw�B'BRnS��a�e%�|x����EҦIM�["Q�(���U<�?_4�z��������)�����s����Rd��F�ն�Q�@��u2HN���;�(�E����t�V+|H��Cw*Tt#�a������e������>�=?�|t�Qk2I� ���w@>:8�A�M���.r�関�VW�q1�0��cup����;�1��Q��ą��"��$�><�Q��2^m
�M�������Af�	%U���Et��@����� kS�=��P՜��a+ہUH>)�<3���2�:!�ʍY��oí�ign�%+��*�X4w�X}=��)��G��ͦKR���N�BK��'ɫ���B���aB󀤿����џc�k���x�O�;m?7y��m�*y�����ʐ�V�&[p�;�����4Y&A|�`h�D�%�ET8��3K���U�����o��IVVY�RCh�f�F�8�U�+FR����v,U��P���=�ja\�����II�Շ �t���@��~��`�R�+M{5ө���F2�1T����OH1��K����6D'��$����ͧ�/�}�/7�zo� �#a�(�ϖ���n���r���+Џ��Ӭ05�T�N�ۍx԰�l���B�������b~�.�_^�d-H����׈;�/����y7� �7������>4^.�T&'2�U"嫼�T,��FbH6�	�����9�p��Z� �_��*�^W���}�M���v��c9g͘��/�>�-4�o�y��|��`��HKp��SΈr�"�֏����|ע���(�.[eAd�k0��
�!�T)F���/�ݤ<O�q��0_Yg�����-Y���A�,z�lh�=4�i���w��d���GĞmPB�`��D����R�%���=���o^4�;R�� ��pl���ʷwWg��n�N
��ss��b�Hvv eK��/c�I��"��T����ͦe�,I�9D�@y\9��p�H8O���^G��i�H�IT�ҿ������T�F~��M�d�N �-��'N�I�V�S�u�����o�\�a��ʨ��P᩟	�;���5�4M�i��q��Zϫ�X��틛N)�n~��l�Ji���TaF���5�~���g��25�"�]Z��={��L}�mm