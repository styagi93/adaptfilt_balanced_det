// CIC_mux_probe.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module CIC_mux_probe (
		input  wire [15:0] probe,  //  probes.probe
		output wire [0:0]  source  // sources.source
	);

	altsource_probe #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (16),
		.source_width            (1),
		.source_initial_value    ("0"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.source     (source), // sources.source
		.probe      (probe),  //  probes.probe
		.source_ena (1'b1)    // (terminated)
	);

endmodule
