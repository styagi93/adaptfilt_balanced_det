// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rTLPlFcmpSP40bp/AQVRde/kOqzf378gbws15OOlMf9DyRyhB9SUUmHUf9jEoAVW
OAwcbmIvY1sSjM31FTyghoU+uph9mpMtKegwjCmzjriZ3jzQ/Fpv2x6IIPQBdG3I
J0inWknuar6wRQnyoeKx/fTejDPn64QFUgorE/XumyM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17376)
xN8xC03wSjv1oyr/z1OrvbR7AILi7+ufnkNLsY1R0Dhq3Z5NFJzwO4gj3f0pPkEv
Ukk8N961R6ds58k5DwjED996WVmHSB+gPi8VXkiVirEg0PFHmHx89Cf6r5hwgO+7
7v7WQbWTBhiK7SG9aH13Ee3WCF/iq+I26jU4IsU1gUKfa8jiGMw1LBbzpy/JxwvL
We9CtwKOsNjLpI5VGIPpJTC0vReJAoG1k9FbOObXGuh36GjcTnHVhuIahQvKzhsk
OS76OSNzLMzBdUd9KudhOYlonRC1b9qdj3rUzHAavs3C2K/Fhr+Et798181rmaZv
X7nw9CIfwQPZkzzElIHEiAe2HjDXDFOSpDHudefBNOJ03WqEi0+VXVU26dl4jEnv
B/rhIrBndD2kru/Zr/oSrjvb2J07/9hfWfskx7gKbC0oUpAzHHs2xFl5dH6VE7DS
ZhOKMQuFafI+JymqNTuhBuBdxi8FQx2aYuL7fhA2CnQsLS1Apna+hvMUHnRQxS7L
z0rZCPb5rtRIDBhDr9CqSwXTWtBmWomVrPZ/qrei9bwMTJUuohDyA8FOlZt4DXd+
ACJ8CwmNizPp+aj9ReL54Wze6Yd07tBLedblZJ6qtmrMJMjH5OTZn03FLTxv6VVL
15GkstKCegV3dQuIm3U+QDGRxkDlcfdFwutzBhRRT8WCHghMT/wFZfeG7Zus3PIR
NOodpuOUhfxqmgX6thVt+nGnDeYmtdpBbls4VRp+Xzgunoi76D6QsXmCw09aNmaG
R0pD1+XPBKCcUrfQAVmaIL0pR3ZfiyNmRGarSVfgQF3wL2gPz2f+6Wwxb/7rCF0F
mF2IQ+LYKS62ojZ27GQFM6WJWPmMWggurOluab91KFLJFCgbmsYC4RcQi7Y7K5CH
5A7oFhQggpAC3PzJQzJA7f/UdNaZEqXKgoY7k3VU/Cj/eW7U6fh8gEXIaYGD0wGW
0OwER4TWIAF6bNnf6/m0rPdsMxtGBGlkNelU+ZK27lw08QTrZRBJHdaYYcwgbkhT
JslQHXNEJn07TxQE+Lrqg+yMcNXaIGrUJdfNquY7nlGSKK6OPH9D5ag5/bV2elaz
UGWnmJcYBeUPZGfEjEJxPLKP9ZWp065HcVzwLGYZeO+GcjEveCfXp5pN/g7GCXlo
CB2Qo6rtF05zPZ64qKqvdJuLEQOufyB2MsjkuYEktWX3SnnVeB2/aRd/jUh2YCc8
TXWW45gccRA3aAHzFb4gLhFTm7Z+3K+vVK6FN8AJQyw7g/XjvizLSGeo4po17Aom
pSWo+F6zvgABHcqNJN49FyCM5h/wsyKufQIyYX8rVmrfSOJhG0N6nQJX4RF/5i5J
LB5BvlodkcDGvKR88/RSzXDYDJzak3PvMqcNA0yiAlkPBh9ZuHxDiecz9OkvrnaO
wcxMrUgdupCzeB4KYf+ys2bTOqBK304YKLj/RP1jrBxoVan7B2d2KyfhwEGpmGJZ
08WJqsVhxlVJTRrqWxVz1W2kJTTuIPwfx0dLh+qaFX+hgaQOfb5M9OcvzFHXEffT
KdNk69d56Ppp1Nopo1UQRHe6l7Qo71v8MZF6EHzdiry8gbZy/jkXiqkUSnqJFDRO
j2uGtZe3SaHhLzZeFTkqCCDB/PjvKtqDnJNiZMEu83rZ2NFJcmZoTgfv3Hy4N6AJ
qXDHfM7Ap3HxbYkibM6SpvrX1d8Qi1MnCezgYIlR724clF3CTH5TSDBrbfk2idhR
GY5qJrUpQxPCl66q8hrXivbwl02yPV4/tckB4z7idHV/YF5hDXxi9CL1dpLckNpV
h9sBvIWUwU8aRODtUgK1JMrryKEcSyPfS9Wd0aMEiTUYuiLYRqrPRofjAgFSVHZP
0ZKkEX1FWH4m8DrPKlhWMrk/JRPo13+w4PR332WfZsqqTvqWxC9ffsUGgBO2QvD9
JoQkW7IiwK1kY0/BIiYdlCledKuyuoCUEwRZ7XsAm0InNnBfkzqUEZ3CZ0NuRhob
2ZR0pZTo7AQPYI2ZVkBIpqTlrwng9pN+I3HTyMzV17lAVGBVZ3yZDiisEI9S1Ih7
EGBEU/zgUqBhewTYHO+I/KFvbwvypYwzIjZx8sSe6N2F9Yt8jH0sUchLAirdEvpG
fnueyBihPl+jLI0xyTygeljyUEScJ1tji188N17Y774IAUtQ9x0TCiMkPxhMMswk
8V2Ddc2GMflFyiZFCy8ziTSLRt2eCpBoXwiWDd6vZY8dnMJsZbpZ04bO0kCyvjes
mji7CZY/BcKfhbbXkvVTpf+XmRMtD66UIjdbUmkQqjkn0mcOoUda2k4J5K554BEt
50mtb/1ilzcbstDIO1pQXMtos4E0vHVKFSqzwT9noZkSMvHUTo1rPQgyo+ldMWCg
4UajbedRlPWG0yYL841Jj9uZXxdmnxLLkJQVQLPw+eIGNwrDWB/mQebsgqqH2nTB
J0F+CKpd0eUVjSOVGxbKYkSeLRF7HRtW7h7OAXUFPz8hnG531Q8W/j9SJgN0luEU
xwFnDeZiCyQqelEFgKe5Ok47+bblllbVd9Gvq6qq141U0d4Fw+AaYP7uHZUir3e9
RFy0cXX+12/hwrTCbOeDFgVT1ID07H4Ql9l7hzOlJaA18u3qWdRvMYZASPmeYGGC
fZKdRhaPAC9gwDa5rSBH7Rp4+qpdCxPwqk5ZtblI2YDZ3FKwqjF26K243yyj6oRo
ue+dTqS7sfZWe15A5z6BuZHsYTdICEi5f7edjEmdwwetI5gJTFMm6VaJHExl6Lf0
CUG+Wu2R5MmVla6jU3SfISa2XDaD+8Hdjy7LxmoiLGtTOcHxp9yLWorUNST//sUz
LaRCUeNlsggGFh/x8EVSPE/bmCnjxEzYnhOMdINvjwYHASXHX7akKAmrBl/RJa1A
tZH+gDjIoBdzoYoMFVlXA7JeyYWtYAeQNydEFrczRoYh3j+3zrcuSSiM71ucsVzX
FTtaLb2/V9OK7efYERlMQoXR5wfJfV5n11J24gre58zCDibTWxE50eFaLbED7eRL
1hqKjoN98Y62GG8ULQXKhpuE7ysdyYDI3Qi5W8qnB1HicvKzRhBqLfjk5qjpnuSa
1FF76xEPb/bTaRxSC2Eeo+eAkGMSQw1bzCBqPF44+fKaI+sSwFSAyJbxWQqeItdp
KbtzGRcDmX08P/OFJGOLk/EXmbBUliN9v97QIEWjaGOn1qjvYvvSJ+4UrxzCpLqp
utAFxEDXfKd0SawRjKZnLGefeCSbSPnd1NtGGau4Rm9B9YX3vBkjiwhcd2Vhd4db
ROniBf4CZq3O5dHx7hkfK+psoi3BG6C7dxj7IGtH3A78CdXO3b5aszKzTXvh/SlO
M84JDJVHEjreCuzmGgKBHlLXciFcc2bwz1dWQMO3kLpUEYpBDnTsai21jThQ8WWd
qanIAfLpnRqv6FrY1Jt1lIhyuP7XsQW/yMNR9dMMsMqUyWV7NphCMuxJg4HbKloU
95oUk1D74fqz9NMY9eFI6BXEk+5L3bQ9QQXAiqpAGNbozjVoX+2Otiqz4+tw9HM+
33hT3xduXWqlAXVgWVc12senMEv7gEPachjiLTJisqR3TIBsjWr0V72QhNsXRZZZ
GBA+0Ec84XovyqQA4B/4f1IQIxNHdE6oSwvVbh5HzHXE+rvEwgkG6a+thGD1WFLQ
5niQ6xjsFjJQB0haY7sC0VFyaLe3eL4Xw6YA5gxb3crb3O14rdNqiIVcEETMaGks
aCSt9hMWiIaytUNIjMhyXQ0dacjRMjg10RsDuAV9uuEVkiza6uATYXl/A++4YI0J
+xbwXz5vW9pzPhxWR36PAR/NIrKzRB/sfcJ6Rvvjdt0g0lmnNDxSj+OQDbCqChw8
JBN2SwJ8xWK3KpKZvxTjZh10ewnqT9+FLrqTwOxROdyzZxljmAHi9Q9sSBUY3lXP
bIfDG/m6B62iDB5f1o7s9oXs/RDrGURG5y7Cga1ZqWjhIPBLSEvmWQHTbfciQ/iX
xAETgVMWzOwun3+qn3bnpxwIsEkiEzvG4OMsbgP9HNbTcWB/FOGMABJ9N+hXve6J
kxaJ125sIFuM5EhnTIEkG+2CB/jmNxG5cFBIBOBHELqM6fDHOhliJzIVtlH0WFqT
0e26dFAyNsSsuFXym+aIzTSELGhDWnDLZGehKWLdFviQchioArgWgj1cqgRJU7EW
TE2XQOin1aV1/P8zk61yp78GWKI6/UFY+mAsNMlSUThP3c7gLfUFGtwXqHZGn+Jy
+2FZQYf3aZyS50fMNQmzNC/s6OBjQm06uTAnFvHtMnK9m9As7CajLHfCa0QPOksa
rMJEXjJmNDyz8zUrUh+nLxjp94emyl0JXT/eTQ8Xrd0cjB7elmUPEbY+eZt3DdH5
GrFELieXLaq2j+tWXH00Ix+QuUSSY79/wSSXJFwuwhoQ0kKocNcC8WzwHVDx/JqH
uuqQoEcYvxq/Zeq12JZpzFV9Xmmgyi4oXj1wxqRUYeGtuGJR3vgOncOUgP6Idfs6
/WOadp/RiNo2uLPSkjGYfl8EShy6O30otwDk7sYgKpiylzPaXYrZCjXnPnyq90Nw
CmpSc/fz6j+D/nGW4LZ7LtsAXqaljmP5+Jq3wPzBVB0W5/eh/bSRjt/DzCLunoNo
zg6UadPGIPx17Cy9grNywqto4GhryHhZhRT83tkjWFhDLlBBDr+eFevy/KFJpUyb
76W4kDKy990DdfwewfMLQLQIRQYwopuPhNvmTf3VaeCLMLu68vGo8WQuUdryFlsb
gu4QDaq0tqTgegQiwNuRqp9NxvPWCD6oP6G+L78HxxnPorWYi5UFwkff4Y/HLDKx
ll+thb3fVrJS0kCwDtkE8i/4IPec1MUdS5zLq4Ay2pZFgftKLS5VY0G/gsHkio7m
cJ0M0aOyfV0jtldEZNBrEXIBUSrrb4S3RWrqC3U49WIz6dH1wjAeFFf5DpfMgxzA
AkUS8DsIoGOMLLWXMB+kIVkrsryVBk5sk/Y4Po2P336SzvucRn4hJpR1USqBYxNJ
QJ56X+eUyP/Mu+3LelikYYCKRl+zKUscCxsc12tBJjIvS/D6ZJ3Z6c08JB/mC9rj
MGEMIcW62AAKt0j2WmfGnbdPOima+v4drGF5BQS7lc3OYesDg4q7JlZhV448dSBE
+0Xb7Plrfb6BzQY41q2fN5n5rfj+V6FbdT47N6AOm70EqLSvo7AaX63paRv0dbME
1xn1oTnyqY7ky+n94nJzHbtqu3kFqMSuwzr/pNCTQd5uL/XOuiAVE1u7B5AY8xas
IwymfHli3JJrYlocMZx20qlSLuR7daxPuMdABTfEKSZ3XcMLPge+302PPoTS9hKt
mOtVGnp9R//33gfMDAji6EsQGFErXTtUvZlu1htfghXZ2+kqrhi89mlVvoX/QIA9
C0qw9fLQPAzv90Wf4a6EW/uW+dONqWH/Yxr6SmdlW0Op3ar2jsUvvrjy59I1xe3P
Y4IoOv8JNELAxRf1y+BjTvhKgP9xHPD0AcYqisZsF0xFbPFp4FvNHihZyWHfJnyO
pOjFKNstG8n/NNKmUcieLXS6irvXQGCVOKwGNdnI+G+1CHCTe/OKlOa2lQsca3xw
Qd1kpa/RbH+3QkZLotIfqsFGVRCxvhbgwdUCU8Nar8dBwqn9K+QSUgNSGlROZ0Bg
YEUvt47Wz4E997sGwV+eS2kDrtHr7HH9em9/8SFq03xOyPwwf/gnTMXsXwnyLG3O
MRftgZq1y3swADn6osQrUjxZ4oFHkO4tEszI5idkm69rniHT2RVO8qS9Q2yr/uBD
eG3C1k8qJ+pBdEBzgXsbthYYZ/LmIiq3URnQI7Ve83AQOL7Ekuf65/co3s/R2po2
1NCJ3vJ5XNVa+iya72uLC8/p6CVqtKhiA7vbgYAibMstJw83MbqiUSSosFOMijaX
G1HuTwfzmAv5bdR+mGhYyWmrN1V010wAigdvhIGy0zCUoAR+65D5G5ChLVU1cXku
AB8Q5xFnmIcuucFYsKV0VOhbgKNs5SGdlL8abme2A7cOWV2tyOw1oTXO/WXTLBvr
f7rX/NE8vlf25jHTcNpdMMBas25wMAg4wQ+RYlmNYIdr/Cl6tOgOfYTAl7m1sS9M
2DYYOY3NscgDkhFfdrb+CNGuzFYuMtTnC/cdlD7ufzgAZRQOzJ8afiDk5v3n2HY5
jcSiv2R0s6PdjQeEBcTWnrNxUFjY7HVwG6HPB5VlDvkBFvLBfgX1vxpjeGBJRr2q
wxAYIoJQi0SEpR7slenGxna9nHVAXXJWY2OtHaoMAwCaG1pe9DDyBIOLviil+rZb
Cl0PNl4HeQcpknS1Msohaas+IrZUUssxCbAQHZDIcyVKdOg1yeaIo+iClNZZFwZz
eBVBlKa2kA3qHULGSY70u0K7vvCUNdvEiobOe6ro7MNUu7KIk5nTMkS1aqRhY33k
54/Ip7Pt6F/lbdfl+1agltD40N7U0C1aetV+O9BKIefQD+Ar/T7/y+TvapUoV8Ji
n7++bt8CUaHgW61KRRTxI8oGTHpN0LoKuVzcx3MRo+VT1FS3ehmsyXjHcG8vJd9n
jVTbU2aTmdkEup65svl1bySu/PosUGna1XdMKvx2RxRlCgDWK5qknYaVD6fD6C6W
WsUffsbcWdCYnDr9UPU+Uys/veK2NSXP4b32AhpLqLgeCxPkYCunxH1FtztaBbHZ
DWJxvZIhMS/xaOTLUGiYZHcayvju9hmd05fgyejaCJ8JP1plFNXcok7IHiblNjlU
zZ//Vm6dkppBqy2AYAN+JB4akrnAW+W5wVCPpCKY8zgExwKzf3P7qH+mptv+D5mO
X3+RkldXX1Acg5G2HXxSbQuTBLVed+u+lT5Ll4W0P59q4lELAtwGVHUxkI2Q/e1T
IWHcGk0J6pylXThTQV2gp3LOXDUxxCADIfKM8j0eEhW9D7umEaQ+4z6Dvu5HZisR
ilrnEPfieLGYuIXNRxJ/MhoU1/PxReS5Le/0kxKTAmF9/2DAYdRmmqsTZFSd5+Wu
JOm47Xow82jREJKqMGhX9/OmXe7fF3o8PIymG7Id2v0f72RjOazUKGu8QdJcQ9R5
cbGrq8xqHXbMa4hPYml3QUu08vQvXgE2me2sZZTutr5998qDWoaL6GTkRCM1nTpW
CpFtJO/4wkI5E0sG+bqPhDgwvjO1DDUVB9eGEKOrV/dNzDBh6EftYB82lG4V+McV
bLokQ6WZpXInJwRUripzwiu5VGzpzevffZw4XGjTT63wVSGEHZFFGXdYiteAWody
JaLtUWRcHx4p7t5PoOUiX2UqXLgOyXtmQiCvwQZRaNtvLcVxU3KZax5iFGz3NYTC
ltFwqrOG3xV7DQXY2QvpmBCYRJQmlDyuWNXHTrk+BNUBj8sndhi6KvZvpRCusqkA
xjtcxdT8no4Wz0s6WjEC45qKj2nYkKLjpAMz+/v73NZS2Pq9qQisq+I3iFWf9yk0
h+1MwgKswFFpk1AnsHlxzlndLss4RmygKMb81uBHR6xyve5/ikm5601IbKMHsrLj
an7RLiddcxtpRM4GX0NZVZlrbAmTXk2dqkc/hChflbQPPVoKRpJ++T0UFo1rsc08
eQhFtNGI83mKJEQBYCLEW/Iow9ChWWbRIMorluoUI69fnpi7bovcDiel7o0MEqo7
xvAbGFfyFrFYgh2UhJShEl04pqNPib5qkROibP1L5tXuSZJfVJy0jZYn7B/IFfjV
XlB9LdJFJ4Rmo/EJq6jfFiAfvBUCs+sLmfk7zEHk2m1VHzvl7o0CyuyyScJNpa1H
gaK6/EaLDQ8vpc5HdMLWwEIs4ZRQH26hpYBHK6shcQRU9rA2Czk1N+6GDZQfBcTE
naajfBCGgnmdvY683t2uS23is9yEbun95MNiy0HoCETZZpyigUfOO3rTKKgXqk8T
/Nrd/RpkknV6vKlH3mQ04kbod3q7sYqt2rI6G5+p+LkYoJee7p+ucSFIEbU42v4E
2YerjB+YOzhTTX8l3qCGsDFGPp2yyGeQPZfhXlPEu9fZyhEmTbp2Yud27G8oq+5g
ud0yDhl7Oae2cMhMPBzDFga0T5W8fsqgdWZWz+2lIU8IPbdtduAPU8kDgguiie4T
6QY2S53pi94mRSH6YnyB5ZnyeTY8Tf2joFvGSjvpZMiVqVJYrJTBiDVJilwzc1AI
lH6Krr5/yFGWhE0w4eB377BFjqR3tzwPAhdM792tlWCBjwow9mB7hsSvOXmqS7lg
tocx2pK2V2uPWCwHxGtK1DvUoQj8/4eoKKRlHz6duZbvOI+BGvX+hg8Iq/wn3K14
1+5K+huwXI3Wp7QhjiuJOrbXpBXT3DXG3dShtL6RBF1ziRHKPv2ylAguR065jQaK
bkfXgKHfVvt3Lx+f7tg5wj58qSrwPDkseGDAVOx+hUjaGMZR5irbq7eeBOGQ0QsO
Z5cszmvmWb85h0kU0vhqi3f2mH1OQQHp/+uSzYXosuAFfrGW6flJCfzMozVa2PLL
BMnouOAEdrC6VwsA6FgljKeWFf+DRkh56alsroRpvbsyeRkZ9fTmYYbDAii1XEal
MtfVFXiTbJ5fyiE2Fwcdn23/sEmtF/vSe4iJUBr8WV8Ji92N0yIIOHWctxMUf9ao
YVMfQyfKR/NEe2seV2HJZWBi87NA8+mFrozidrpkxA6RDRV7F1A6aV9kCsNQfvik
OIfNDvbHZwPOcQBYXn2OA3QiI6/QKhBn7ZmEYMsuFqYnSv3WfBE7yRWhE9dzX80q
ICaf2w2Rz/ofkdoVrQ0udAKIu326DkDQTdUZKcdSSI3scSR62I68phEWSiwAmmzd
z01iWCf/q1+m6bEHgK15kJPjxFrtfjyLslbhyXnd5lpmtfIH5l94DPynZtvmRVyU
OPsM7np6KsDrazgIDPl+8KgY+DvU3kkhSYPazkWAbcSYVj0ni7NINsIc3Q5XKPTq
rctaDe2TCSCzlsP8/ZqH1+K8jN5kKFPhZ9ujjL1xayAxMmKzxfIcfZMz84j1Xumv
1gvifhJhpRcYs7K1qv6nNG4Uj2K+8eF8bnI/Ex/kfJ+YpX3VOdX8bMrcGcp9ipzx
94cA1cisFiQJJpOa6hpREgvfBwsEiktkfheK6kjcUbxPUppKGDgbtrvbrLZTMtwi
WtSyVY7A3ryWEUX01zIxvnV5N/4bLj24K7yPwPhvTArT7kKjru676GFJTzv1RK8j
4TzXC38eLXzTQ//Dhkm0BaF8Gy1GzpmtsvUNjtyvUbOX4t+3AEuXFgHwgu/0UBTS
0I2qqCecWO9rzzA13JcyfZdGPlcQ9d29HMZAZkJIIxiDTCq/ezQvmnqF9jbOLIP/
wdLWRG0XiYLmbjQq3+AFVmn/EbY95OtSohBTXBkAL0MWeT01/sKZihtA7FHicQJE
XS18AOnu56ZyBzGeSdE5iEycSbZRI5yS6yG6/IT03eocJyAlcU4OsverMsg2p3jx
SGUJnSd6OVx6nm3y0kFJTs+qb19tnmsF77watL5HHBDpUctxk/8hSjUUA3k3gXq6
drGZMSxhT2jrGp4Ri0RtwVrhaynX3JTsuWdYHe+qv128OLNLXxqzqVj/R+GB/9ks
881XobWdrDIJNsx5ziNnDHohzCmlFf5kXhoipP5UUIbFoNYRtNFw53viHvJbTZFv
B9lWGbk6iiRP/kVfsf35j3o+MfIP/KCWoXLFRbxO7JC4F4ZFAeKMi7gv+MoQ8w3q
8/165h/34VO+2G1wYXQX8T3F2VDZUSQcxbp6vr/cz9FVmxevbWkLoEW+U/+tlrjr
p7r2Ba5DpAlLZQ36S43p9P5ViSjxqqKRRk/wW5NAzsUe5vZWWSL91yjVQL2tB7d9
xidR5azQpdH2NMcJW0rk/l/xSp/MGtYKs/csRsST1kTLQZVcKnU1ei4JdVB/FXlr
nHUIqFNRpVtgmc2LWFMX/loKYnGNb3gXn007nibMG7wO57lwNqdcKpbo4zTe4V91
/cvop4tC8DAfDzSHQMC5JDfT7qwt9m89bxw3RMDrAsgKkLcdxYllTK4NzqnJp9FM
U0hlyj+ErcutcI1PAGdwWOgzT2eKT8CUhoiPEbBjXixiUpigBq8TIJQAMNd+tMgK
v0qELgK7jQsZd0mG2ch/kv6Ikl2yM1TCCbjd0mE8BTaOJTpkR/EWtbEX0AydQWnc
mgh0UxZL+QRkfGTJDGI496pDILde8cKcnUaL/Yz9nP9uda/i2l4bCu0LdSJDxDVY
0NhWVTMnWj/4kJN616ky395neD4RlKzDEKa2lMM6ayy+X4Ww76nkB3THZZtB5GpZ
snhQuDyYsSt0viyY0eWotwEsmsksswRWdgZbEza+VQBE1TlrFqdo70kcrcmlinyM
F44z85PYQrrc3kLF0qg00KZJ0VKPNoCRPOeuQwKnEvGZ/LqhrQZXq2tTux5Sd31b
BGIWF1dORtN9qMAHnU2tDnbJ99O03P2q7HSRotEtA/S3cQi6+iRq6bbwtEgtRiq6
4YStqqWyaWW9lptahME6cyKfEWfBct6423LeC+uU4/mXcILnNhOVt3zicveAWZ1/
SVvk8vO0FzcN2NIlt15dGn+/ojPkXLjJhyFhUExPQldcgTb5/sskWs26LDNEcrSb
KoqbmxLR6ajLI74RGjblHvYdWv2VzEW1n68q9DBeeZ/hMbmfvHSUzwV2SWGG8sRY
K71zkfpX/NTwPLSZ2ASaCTtq6CR1jYRako9y3996VUv5z1FN/WOv+3iQC1CPHejq
0q2fkJge2506pY3QKjxeY1RP71r2YqstoRASc8xc9t9w1BOgtWZiXIlObo+oqmYl
l3pb2cb1gZ067bOcod4cZIUzmo+2Yd7TILuMs07taIU7pCOqEmTOTzqDmLLEZTDd
QNeKsIKZCGBFWkEmI+W/XSc3ZlFSPsEHvcxItcS6wQ5l+a1DZNcTyN/5KsGoPH+e
UoiHr+/7JWXIofyNEYGz08CFKH3Q8DGBVIk1MbOIZmKBdJRQD1bZeUgOc6W3a+fz
u/qvJf8ffQHRso2ljmsPJViMyxs3YOatxQKbPyE9u4boxMFQcerB1UUw5DEhVC49
7mJBnLo3iSbHFnAGeffdLh58Fwu+avoEZ9o3K1lLeXPLa6T6RRE1sE+thYHgQcwX
cyId+GrhFPOoSpe1XJTWBB+GNxqosaEh32j0pxbpxH5d1uiMFNRsRGiVXumBd7GC
GFxn1smvxDNIX9wrDem7qyBDEgALJxyGmWpuDeG9kripq1sJbczxCPxN9Q/7exaU
o1Giv7yf7v2w8X0YugcfYGJvy5QgiLoC4P3FJ5OoOcSKaWxwcsVSWDwfYyEawd9M
P/GI1h91bszjiscmNWpWgGJQ7QiajMX6Q8wHDFO4yzn6qT0yr9xS2ABxNruO+x3+
ChYw4JwsgukcOFJbwiZlz7OAH819z+4vH4jX6Z9wA0c+WpprbokgpFhFEDR0KMbH
PH7WBWZa3/6QinQWMlX8tnV8nI6nuYl6sjXKWG9sLNOS+y+g0tZK4y9+mi+apXmw
qv2JmbUgys4J2KnLs8amXSEqmRL6yUKvzcT/R8bZk20VXrSkjgAOW+fayB9KJ3nH
21pBrnQpXduKSrrz6LFSlQWcDOvs4rcNqgsu6VGkWm1zcDgp0zDIpMjkAe7mNnRz
SuQmRBQAyv4+8qRnQ5j+x8jyuOVdo+AJ8BhG4sX4vjoksKt5HT3t3BtN8+vMLuqp
Lg45f7Q4boF4SGDjXQR8P9Xevv2apeOpnoQQ9fNTrMRl4knfmhGR8BpHmP4pDwit
0El700TAigObxj0ljC5hqyYv5UsohoLuSJs4iBpR5qP8crZq5shIVSskhIJLdZaH
00DB5cYbj2TQIcS8/mYT+fSGTHk49xdasDQRmR5SRFh3Bt1kvJBnXlGjGPFUyhOK
6jXVcb6bbGHV1BRm2XuxJakW/DLDOBN5FUyfAgwGSGsDD3ns1tq8KwD/bCbbWpeb
oxQWsglGisY1YXp+JgYfNvA0ac91oNBHMoIHPYhcenjRkfRqCZbFK8ib3bAD/P3N
almIbwt2QOuAqmD8c4JjDpATDhQuRBiEAzYUVfX90L11ko3YAYnKYvhSz7Sp5jNd
qxbnzWPE6m+X24zvE3nDzAblYGGBlYsEbrTphpvWd02yh/d6wDrXyJtse9/wz3fR
kJUavQJo1TOojXovA1SZPg4Lp246y1coPhcIiORsOdFn2DDf1+j5lhgZqbkILW5+
RRg0KmzSW/EmPsGMjqOi69blEbJKqMqnzK65VO7m3gJBAqsRX/LxBzhW3fVAWoyN
K5y2zR47yqS10nMrWsjcKwzgB4FlxfXm0rGtN6SvHRT5KWnksvpTbVLXBCi/GLNQ
7KN8VfHBbdXl6WAYX7hFhpBsB+y2C8HqE1wntBdRi2ny5wQcrEUXlEZ4crSzUa3U
hUcFf2bCqhCjS+BMLSlf8l4mI6dNof+T62Nb9UFUMifxw+QZ1zMKWzw/DQrdckS2
uPa5B7XjhjNJfJ4L4iXO1oPuKHTXMIYHCtmO9n/625aXKGrC2vZ2m7G5vj4t8YKy
hhCInJeHuDp3LwidpJ1XCHd/Sl+MYsBoz4tB2DKiwawWMw0jnYyUURnbRkzbQxfH
4wTcMsaf5cW+z9t0rIJ8yE38lgo4Y01hsPFkX1QvSE4ZQCXCDeAtsvBAyyFSc9pp
PCMfdxZ1i0yfbPDGCYWy6Ik9RJVT96gM6taDRmB1drxHJXY6HtYDu3b79KLRejpx
qrrfsicuqh2IWQCKpUKAt8aL2gQgJkoH0EEn354mBqhC2EQ1PcjVpXiN1FYO/AW7
heCwwpY6+W45QmcBZ9x+ze7r+EUNh1kJ6sxF7+alxfu/e2CQ3yxpR8vmwt2BCRFy
8tVsWSdvh4R3LizzGI/JPcx8b1jkkRI5Blsg63b/B1n6HKtbF2CCFyJGdRr9TLQj
bp9hf2mQbq30zTezNeTi08hVwLPVhQyRX7dUEWnGiA/jWZkN5LFEjKQCeSI/Zlj3
Q0JKNs/dnqJbglEVzjBTX0/JnBHSWrGBCMQxlRUDJ6EhcCgJjry90wBBgGp3ykNP
u6lz8juifYVSzw4dEeuj+G+dr0iqsieROPY3zSNq3ETLoJkmNeJ0OnpkkY70J5VG
omMayqOYA9mbv0xwuQmQK1mioiZcM/++T/r+L2nfFJ6X/08wC1SDhc4nt4Y/bAnW
5jobEiFGy0K+Wco4i0P7AHADpOd0V2v5rsMpR2tFvFjVTbyWw3HHj4V6e/RJyct+
QdlP7F4QSvHydZAaCqXlciglt3jIn/FchzFV9A9GSRyeIhPXKWb47Mj0KWHB4K5D
WHSENzmLbPJTCktv4UZN94By71lJrIzcW0ZZwc/IJmeCcUBKfrKw8Hxiti104xoj
14wdXgdEQ4AYCaD0muHckKI1XMtUuqIqIIgzajoJfkIGi1Q2S+bvSel0+WG4CaUc
OjmGk8Dkh3dCoD6ViJOEKCN2rXPcbz8sSdhGOZoy7tZYSmRdq4f5NjYL8X0xj1IU
1/devLzOysg6bDIhzvzXlg/vJNw1YWBH1BHCbLdrEehdKEmrqTOQftd9ghL4qOnW
VsxrMMp6RxT4tHTLfmPNCsgJCBU5pUsyQiK3NT1UPq5BpygnhVZs/pwBl4O548cE
JwA0cPXiH6Km/6+CINGiwN5dy0po1ZGEpgr+9ZyIucxmXUMcyBQ5vL7VujRojnRc
j/NqXMNcllaKC6/DiPuBMKUJv36rKmWhRi63M7ZDSy00QuldFH5NAU7Rr/rgRnNV
vnxOuO4s6cliXed2Di8+Ll2e0IJ8wEcouj8niIX3tTxLx5OnSs6nr5WuI3qfFltc
JsnKmfB0aaNdlUvCB52pC5uKJbggzbjwZTPMwhjqMDMSmAlCt126toTifQYg2bIZ
0Skp6/fr6LebzhzWt8PL779lUhiWtn2he/vy3x8cAm1yyautl48f937XbCHvmiko
kZP3wu9iBnwLIry8HTqmzAf+n3S7HjzdkCta/68Dx+9OFjANOUSxBxCNOuY5swD+
2ZdxRNheV5Zi+XU76ugkI5EqfmecUABeGXGgwDtb9WHAYLAUjZ3/fLKRayxAiuiV
97FF7RwwggDpp5uNTZZZsRGON7xXZd6rPP0K7giYgDTANGIxOftD965eiBeqGAzV
AbFh4HcXbqMFy78ZoH1ZiYHcQBmEFaiPCOeOtQRuy3t1DasEFRgBYwO+bEl5Rnpz
CqL5i/W7+i/y5ncBmh0D0rvJrj3x0sHAuo00nR/PQ2K9ez8a0vButpRe1cdkjL+/
qi3Ws//r8oQ0//JECq/tl1bRfxJvKqBN8D0Nz0Y+p/doJf4cztxp9NhrZjS8Wzno
sg0/CgifSto7UJj1f54SqgTXwgAPv4gqHu0z8GMH2EbRgIsgKa9waylRLDEbI9dz
pqiFq9i7UA3WvDYekgjpVcfUKXMK9PNzuD5gFtLL1FZHaZgFICdTmvvUmcEwxUb9
Eiq1zJAgmvjJKGukzqTSEkwne8JBOvuoQhz8vB5tvd5GmvYFu9jlxUBGX7cDd64b
nkgSPdkTyXloCUSQm7TVuQFVJY190+Vs6qhoxXUxw0Rz2sqy1GWUQW58fUGVWW4y
zwTFAX66WWK1NkoF9COeFTyS66kB+6XYLcXpTtP4CEi3uc/I+UWQ0QkCkp9nY9e6
08TrxXnuGEAHPQ8uKeprv3YShIXaMtMntApdCrSN//SO3p/pZQIirrOFHtELyMSB
fUVJbruK3fw/JwhDHF7SDteuKf5rIzoS8HmqJx0Jr5WqyaHtsjbgRtrvFJvgAbhx
+w9In0vlX8DUciHxwSkGpE7bJ8lA3ANdDHS55P42+pwr0o2vfDRlBBPBKmvDoRUq
EV2ceYeli5YPUbjj6UNmVpGR67Pwc6NA1Fl0YopTGTQihJRcsAZacjPhO+WMYBE8
f85NA+LF+dHCGs7vkXPNY4a8jd0GIHWZxgjFoqB9gFUTYdYqrWEzizRnBus3p6Ek
1OKexXgvwlRFxYjPFx6T9AQr4EQyDNfLkVPOzuyA2w3Qt14kzmhGeLeseIwCFI3z
rL14nNjivVF6wxNgbLlS8iGpTelTauUn91uDNI6vbgt59JdWTlZp7AdpgeF/C/fQ
p7czSu+/QZqp3n7N+zOGqwSN6IuzJLfZkvC30JFWaFXa1mkETwmDmB+Izs/tflG/
WLoaYssmkxqM6JPC7bxo38jczQtNKtfzLSocQxUSaJhUCY8fFJaIXvlZgUZcNNjG
5btQ0RId6BJGIAWhHgsjrhkBH9/ir6QVg90s0CdNpplEmEB7ky8qhKQIZxgAKm7U
mX42nh1SMG6zskZfHOPEjdtbbiwvqLoRUwbgCd98uBHtOr7bIXGR9XYayMpRgu2L
Ys0x4Lo0PyMQBjAMmC5VFeigfli/Li9txHfJb3iI0V+yXilgkzcAjXQEJLwyQUok
+ahtd53sJr0Rg6zdfGkM2fR3NGeQeN4p4CF6U65q8kE4styla6CbwuXsOV1cVImX
585JTYjOUznIldIC5itgVEe2MavjU6Y4kRlhztxidD7i/nTVj+hxHhbBThN89ok9
tHcbLIViX6VwQOFQBGE3yLyBOlDViseWVNKJaVKTlP3Zvt5na9KgAIpMNiYXZ27M
lza8IrH2651yoiTSbZx+617PL+/eazXfZhKvIXpsUfd9OFPyYTZfqiuJjVyHr0pY
KRv2R+4q6VnB+q0E4IUN7xXFJm27P0wJUh7YljdqGb5JzLcFgCzv20O/y9hFs2wc
wGnOCx1tKQ0GU6T4xqaBzcDTRC1GEl34hWWIY8bbBBaALCZbhUaJCiCJIpYWl0Fi
65YrE1ejmHmJSjGhHQcIoOHwoHK8mQrNdkZziwOQDepUvn8StCFQrwrHsvIUNgfc
bl1EM8ccucHX9ckKreaPmab7ob4VjNUg+sYoaO50xV6W6R73iJsJe5i/ukNmp8wN
4GORZeTftJ0+8pMHNoEajURNpJJG/tuLUdCqlnemHqiFBfAL0HmSLUi0wGRxU1Qn
nYLDHS5fXW6XABGvKHNOaGGky/D3Wet5uYkeS25o2/KEGs1ctc2K/hMbNiPuTzvr
qXD7TAWoitbiok3ADNrZEg9/e2iS71GLDj8UlY4XDhynGyVaYPzWMTUFL/kUfVbK
Z/8S+R8juUM0pLGAeBfozSSlmILMvE4gyDFOvY3Z+a0DEmaxZP7ASewM47Ms0igJ
F0M3znOc16tqVbghFqWC6jg0PNwa5+W5qkBXnieEnHXulYrV/jCeLTjusj0TqjQq
3b9AJISj+1iXAMRuzNPuiQBL4m8MquKa5iyxj/oOjbtYS7kN+H0RdbJgtfbEYUGh
XVydbI3ADsA828xmzfu8rqNgxNq35qaqYHEHrJexbwh7Pab0sZtjgVMVmvUkEnID
RQP2yYvv+/3MlJacOM/zF7t3h0NMTywWNna7YXCajZyCSrbDeWeN1rBQK0J91+MK
r66U8jg3rjBcIVfaP8m+fu7Kes0AaA/AwDbHw3GnMXVG2sZHLhzuV22EYnM5GLh9
2xhzBu6kgcjFA24iANpjEqCbuXZHcW2IeVmUUTlX7MP9YaOkC6qnWs6kPxdL+o/C
/UJ4GkPEgVm87QAarzm8QWeiu/bwTeLcA/TmwluSbmM3zSCt0NfgjfNQCm/H9K12
ka+PkRWm12loTAkQO3B56xe7gGOegv/w37wnLrrXespgUxucNE/Hoo6M24GppymR
fffKI8C8SF5x5VuGTA4Yso42EK70VFVkw1efHJJKtiVlSIFYu5C4n4rK85zfTmp9
gFHj174fCM+aYBfrvmAgOCybcLdCxtJbAEK2KbHTF4BTKVyNaUVDhZhtiY2GTxEq
eSzdKZt4wWq1Fl77bC9CnWbhHbbwyLcdiQ//cH0bjCqaVuIyqMi8rXV4IlBSRJSX
6+e1KkyYgF/0VGbf1warmKPBN0p3hzdK0GG1WCiE3hDW3Cnzvgr+N+wDFratTd9A
UAFo2dMTFl2aIyFAM87EkLFVMjwuz+m4AUPRYe6fAW0rRztnlz5q1vh7/QvTfXYN
ogZiZGesUk82vKJENy24RXGvtQMmsDi6CXggtf4EuRju8vv/kyJprQNVwhR+2xxm
Gh4M3WbAyHyoVo2swJe3MfkN4p4Su7WjUqbi/pIaDT/CjuoiEDOhm3qXzfrRzvi6
0kCh9H6inZjlUkBT45VsEh4XhDjPCV94wW+2p7wQpbEZM3g0ISKkH0HEUhgIA26K
7BkCR1MH2ZldQa65FUXssO6EFs3x/TJI234SrsFBgEYS+3JgL5QMJLWJxMbmsny4
zPCe5SLLiKPZ45h1EpcazWamfA9N0jlV9DIz2XjPSJpkJb84vVsDW0CJfiqRhrOp
SjcqzJc3c0c/9pb8ig0EMaxYYnkNC+COKugd4x5+KpEovW6fNfARzdgHEZQIXR9N
OMIV0B+w5h7/V3NZ6LKBb2DfhVJLeTOpFBoguu7NWn51knmgoEywER2nYCH0kCWj
OFIs+JlSD0ttrC6wF0bTsp4Pi8gkQMoynVRb4RgvrJFFo9HSAgivEYwGM4RxH3A5
EktQvQoLVDNNiWLFigxN0F6aSKMzEFreYALUInP1juGI3DuEPg7gdwaT+yr/Vuta
VvUy9bVGEZUvpi5FbcaDZGjT54n36X7NGV4SGYj7DBaQN1ZswvfbqtmsrahgehoN
KTBVVKB26m0rcgU+RIUhIjmPJEQV/stzARiWA0aSpBS2ge5+sB4FdsuuVn6wfchA
etyx2TLbGANpAgLAaElCQtBS+2CCLd/D9Ym3vNp0A0PF9HrTCyih/AhU/R1nQx08
T75kiis2po9jQdyepCylohfBD5kktlCnCUpkl9aNOSr3rKccfKqdAnonxvojGThd
amBsxA61VZc2/msTXqKeDuhuEnvTpNYdGrnCaXGkizTttWd2Vd0uPG80P0j8C/BG
jpXgStZZEDXeNHpqxUSwvbAABv5Z95aN1FNJe+1QuxZtF0Pq9by0lITWz5qt0d/R
OUSPEFqaj6YJlL6KyajXvBPbguQsaYKH6/Z8j6KtrUu5WGuougmynbCGmQBB5XxF
1VQxJQNA/oA+W04o06u6bi9ujP3/iWPvX7szzYSTDCVlXmNlLO9ulNPzzjRT8jc8
bej5G35G4aUP+jqqQktRea1vlE0/q+eZOB8Ze5pDfT19Ip+ZAwsXlplxF5nus72L
VD1uQ5KLrQLRiGJq1tMiGws2RCgt3T3b++eSPRfQxJMCfl0ZzqB8IgbwXJ75ZMo2
1MeWfqLgZfZpcPzF/eSn3dNk3LvSTkcfDVYpDHab27fIM2bvbyASJOzp2YoVYeDM
jOSL7oilb5Vm760NT3pHm8lGiyCpbBDxWn16WryrqLTCGvGfr7pDbLspyjitNHQS
ZvZwc8KBUFHlShKsX9r9efDLrNBSWIw7/+VZhxLt4y8ia0PZm4npkO6X2RTBBwCU
O5hhU9Wv1c+hlCKCEY6JyRD8T4JmbCfsjqJofWdxAyuc5GbavkfzYMMD2anDLmOb
9QSJ749eys1yuKUakRhHHoRST5ymLJzd2seaiBGqC0Bp0WaS2SRr127lVOKiNL8N
A7xg5t0BZHKrpEaZGUP6PqjJF/P2oeJNAiL7tuZ3VDB1uP/rcWXeeWYdchgQG7CU
AzUx5Tr8mFE899e4cn74RzpTXAEbupnWrI2fz1Fpt540363Xd6bSqseZWBww6V1O
kFH40IjkaXI78ZMsu4Bu4sdFJ0wMuqoTTCNVCnNXk8oHxHnF+puVQvk8rCHlueK7
6YkW7YTFSZ3ApqllkvlB0eroIyAZdNr/B9VYZm/+TczsEN3bUUwq9cc8afC8Rn/V
R/2OziYDweRWBom6HMeFCvM6rLxQD9Ddok+Hu4UWGDi5Om2Ti1av7sJAbFlHvQcn
LN1l0jSfKnXddvs/ftdCWmIUFi07Mtm7ILiWgb3iGBx88FF0874JbxzoxmhTbPom
R1eWNcaawRrOJQtClex3qrRpCNAr3vA40PCYBP6UwJmI/Z1k12S0Vge8VPS8Th5p
nIyfIukqp/KKi27idmHy75NOQDeMlOe0AzRtxrlc16iJjwr6BtrKfltCzWQFnqXs
Am12mhGcgHkqv0JhUUqbECFGyNbO/QqiOUT4BgZ10OoPQM/m56PMCu/+gDIy0q6F
5q0Tp+85AJoSkWkfdFweLgD4pQERst4atqwvd2swRluUF6IuUkcr9+HTVJiR6fzS
hEiX38ntugCmnNvXqmin/3mktWJ+scRKDHzz3VAKdj4AUmVsngiZnZZwlmmX9CFE
IVf1iNbOxUWqxB2zVBwnLrhFsIht8S4iOB3CovkCIV+LV6MAcngYKvDKkaRJXP8u
4fIEbkFOQowGqpuR3DOUPT5FgwzF2ZQ9+/VRKkKWN0w9vQrxOpDhlKIv3/oBRKRg
T2/2juj+tTxmnhsX9rtFO29cdJHCI2fFz9mZr1GiP9tKoPY8q6GIIfqSydmXabDs
tAX3J5n7TzNJCOPDGJCAK6d5M3y9jI/UrgZByyaiwMk8JjZrkxXpeRa19Ff8rbif
g2l6Gtq3ZGE5UDwIL0CWuBhnA7aSLpDtZJ+wQAEdfa0IUR5agVDDG+9WkJ8vbcmq
32BALMNrFEKWBUtc1b4kBRTxicRS+XHIWTemJkGIic3QzZh1u3Azj1NFgnfb6ecW
dFfKMHkDhKsvs/T1drGIlXdwEd1I+TjIG0dIL9m+kq4aQ5VRwVutFoxy9uPH0pP8
rIMe9/K+s0wUm6JpyZLjoxMH/NYnPy2fLSP3gUFA9n1D2zHJtqULmjC9F6vKR58X
y/WtZJfhksc3cqhOUcJT5RK7SYIvWRTJElez114OnCYvGP3PJhoVjB21PiDYcbgs
0xmgJC77gd+JqpeTcDcDbTLEqwnHMq8cSSQqeR5DJq4PzBFlWOl/oCPv5zo0d9Ie
qCfc17j4WvYDxKmWqPRHRtrpgzJpN0ZZ+9rBcSSubGGGHzS6EBE0bWsmVoGvf3XM
nppfKS4yEkrpgtZLdxMPoxy1i0T3wT54jGmV1f0thCfINKwqUdnvUjwp4EOfgH7n
XUV7Wd2shI9HDRxSjVSDVQO/S06szyHhQdXbEZxIeMfK7tFNkVhJKl9rH0wlaLxM
ZHVMyH83E48JW9MVFVTeSxaI0ozzi8Q/k54mFbXLhYe4yILQaAfSYUKYUf99zQmP
GfayjxkoQ9hP/8VvyCHE+vejTINX9THNmqNu6tNXvT6TgUDj/YNqMFA7llYSxTI4
2QtXEKW33m8Cc29V8Wqg/tSR6lnUUq2MDnNymLlW/JMPaNH+tCvZDfzpWl5bqkxn
4sGCeG04dzYnnaOArg1L+wmoGpV1C7SD+vrRzwFJodi5VHQTZGXUzjy7Jq0miung
1DM0Xka5RQPhdA8if+QEPkfljQKqvuOPaa8xgSajwKc/cZWoYO8za9/EUZamK1Jk
l+zxQRqr6CssHjCQLH9neBJetuwrhv/Fkfy6Q+073wHLFtXCP7SFq3cJB9YkjvoM
aq2pigMPQLkmYEqkhLIlsfznAptKzrT9n9R3rkleUgeKNVBbNlMiymdO0iNe5XH7
3RRO6hbfwqUE+6HGh+3HKs4e+e154vrrwcMGVKxhS2yWWKw8WUcMnTTbUsdenAua
w/bi1AEplMzwNHFIQJAT8Iz7Fh0JHR3jlDCYL1oXJaIuPXqgvy1CPtg+H7IfBe80
HVwhr3P+nb+CmKZlaae1rgtU/gfoo7erBreT6t6cKGE6tncyE5dHmVMjkrBcYB7l
WmH872VQPPmn4KGMZTqJZ0gcJfEJHh3taaP34JxMHVdQqNwKebxtXZz/0S4gOrff
buLwYjei2v9UvKOkcGZPQDnVSEWIhQNJtLSoDUWqILqPWGlrD67d7sp4CUx9ztAB
usDTLw8KpoT6hpwYjsoX2e9/s/i0wx0G8UKnSBjfnsxyIIFjFQKrORqQctIshrSz
RTZRGqeFO0CmicaS3s6Q3uBpeF7exaWQ/vSNadn0KAcWP4Qy4BuPoUxxGjCc1RAm
y6o254OFK/wZbgF5E8LxDqncIjcj7WT2DjR1s+hM7gDDwUzgnKJDmM2Sf3MyhQ/0
zrbepQhempJqAhIYigrdCcAh2VyF8wK1IuRlIhL776wltBmgBnW9LKicXeFN4/B2
6DzZKOr2N/2LGfN53Utcitqooi/hegNC74PjKRtdRiItoBcAjVm1N/SfLuu+b5t3
e7hYx7vZR5vTj4oXNfSMtubrUnlrrkqoLgn8WWmBq9qy52jkYcfNAdAgUjmc/NN0
M2qYYAzShvYk12W1gG/h5EYFs0IdV4RYzB6963MQAQfaaRLYLM1mVGzb7T065vcI
wxc5/dkrqG3IwPGCgRYnLWUaAoIjaeJDfHdQfFqoJIOmqL22ETdM50lCHsuH0/Ns
o0imJlZwRRJIJ3mrwF/slq9yHVhAZOHy72zxLjVehKvnNZ50vXJBz1ydvFlwRPDh
KZTFcN0nMGKbvrq3Yv7FaZr2+mz7MkHAOVCt/1kuk4fG1/vaP4CAb2HcEqKTliDu
jXnDkz++VTsK1Wvym27XkGGifDZE9Jfk8bzQ4I9WCJJ4WxsbhmZL0bBQyYt7oqSE
wUpQ/9fZIQ5pYlCaVUHyBybPCc6FKGYeWPvI1KddJyqYAAk0yYaMTfRrTwnaZ8Ef
XUIYmShTX0KBjnn6JVjC0LJ7m8y3laBEWMcgLCK3uwYbceL+J8efr1OpK/zKrYPJ
O1yV5ZTsfjcEUCRK59TpfVHUErQdMuaPYF57jctO3m3GVlcM+TJkNs78hUm7q3di
wnSwx7fzimWHj+luF4jQwLqFPluro07QN/kxO3hpmliurNFryzACzn8xBIEBMAaO
T4bvUByUo/3p4lMKuj6I1vRi3ySd54bJLZwKQocLAyYFv5+fParLy+ARi2aXTnYF
LUlUXQYZN/8hbLtsfT+OWT5uRG52C6NnLURXR8pulFK5V+zZkyjH5i6RmqPcNAiU
DWQdFI3akcvTRJBKdBJseZNLiZkpaxaSC2V3Vm3GG9uoWLbSM0JZlKf6vemaF81t
zTHf0IacUL0g+s93BUfKlQZhavpLm38iBoq6Z5X+MqOPqz+9xW/OWnTaezaQVgmB
Pc6ElD7YpdF6Pe9Sf8gUsqLowk/oBWuE27JnffJYNfHAi3obx/GnHzSLZ3AR7CrL
fByLEvU8qMDpc1pIjtMm24OZAM1R0/NnHjAHF7sxPT70S80tfbxPcbGFYm0PzIPv
8kSKno/L9vmTrgMe37Dggdhru6C4HvgZft3KMExnOKSOCIoofB9MX8mXiEwfDWIJ
UmdoSkubrQYcm1k3B2Kk8l4/qFQp+hvFzCXm5llCcKqdpnN6frTiMsA7sB6GGxM4
JMIINUaqvW6ibsoKtpAhAqo5KEqmYj7JKPDk7mkLDNUOSWReVfG82HlI1joulGMq
EJ80SW4rTghDehePu2SGXJ6X8c+r+10gSoNVx9K0EJ1RwjhW3/dAyJqtddSwbtSq
MFf2g4DdlFoUR89gQhw1xR3mI1pKkvWvz20JUPsxBEbHEwkdcTaVlScw1iRf8stn
ZiXbfpehIuNATA5+pJwEfUj0ucrG3VaR4tOl0UODRP435ZxqATPaiaSlUN80qxEU
91+dCoMELQbvqBRbE98a+AFUm8/iVyQKZV8jEpe5P1FCJzAM+FmdI2OS+ceAFpvF
YX0+EbcIVBYG2OCXHmeElepGbxIHYeI4XWyIdTFwqvP/Ac39TaCQ6pwcuaP46+zH
1LZVkXoWOFsPX5ZoszztBlkBCs0RjFbuRvw52CDFHHsGyAwrLvIvv5qC6eOHQ9K5
30IS4K9opSskOa6HhrhvdxIFxUFIOZ5BM2FlR/YXH3O5WL454474EEdS8K1BX2H2
46uj+yxbthflArggUHw39QTIHAxWyNaYTeyqOpV241Qx6Me/Ybd0DsZTvgfqpYlw
bzDhwOcuNyyzDfHoFwhKsuFXrbdxTVDm32+hM3SSmFpDaCX9x8QQt6cPUxIXH18o
1vyOqkAKzOp/r/oG9vEpaKETnuOLiVmjSv+1CCxnnzBSmCDFpxWuLeLO7RuPOaTJ
t+hhYtGere7EW2G+e2x6jkNedE1SjMF5EMwf9On3eCi/J0+wgosJdxEifDtUqZpt
Px8Fjzp7TPvNO9OGtWtj+dNZJGhbZlVGZKIwpo3EyAsu54i/yLftscQms6CDmZr2
TsDJEigcbZ4hsyvewMfJGN3jABjlya6nrhzcMftE9EGfXDrMtBeikJFueaFiQcow
`pragma protect end_protected
