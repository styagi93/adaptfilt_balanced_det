// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
dQasUyOZx0OpOOmyxbV5j12i2SLcbkL7rMtQaYIhDM4hKnUPftnCIbRzoIKSRzcsYkKXukYcDIyW
3KTjXEpYRu2P1a/DU/Iq+jtn5q4hU0ZppDKEyP3t6y/Qya8zwjEeQIUZmoredyXrF0XlLruPEqCB
D0cHnPcJYLkmVw9K9goL5BCclyc+6XtZyo6oXFaE1XSktZC7vZfXBhqp4/qZOt3u6n+H+UauY78g
DO5K6ufG6/JiFXHpHb3JU/P1wxSDjZVwWqh0aHp67B17PjukeCi1inTqfkq/USqvN3SJDWS0eBFM
LgLkHoAqq+R6r4vMbk/rZR2/pWs11GSVJ0WTqw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21216)
/OsjS8udL064+2IPxZSRypdNjTVQ426IUE1DUHGZesbFkaHipZyESGA9qDR5nPqHD0qBz3JorKpZ
n2b10Khsc4Z1NDI8NED8etOKQHvByb5Cv5iZEPgS/DrD3SDYQlphZb1ZBumiTVYIvAGx8SrY4N5n
YQUcKz3qEqxPyzGgmEinaigrQ+4BIb2emQPaLHqISpWlkZ/MV9dj+/s8fZs8Zr01UkZBlDZmb8/S
0ltElEtDyEbfEI7J8ZRKqnYPzCeo3BNG5xoRpE1itH11GxRx+LG63L7hGUYwmBNRzFIMMH3GL0s9
zOXUa0Hi/yQIDCweW2hVRT0iMJedo3R2BxCSy3bF7Yjx0MlsumuM1CZx9wNm09And0wL2KuUCC+J
16cFp4hHzuIYez0ibZPY9bcrbq00mB4gN+oN0+hn36fTUm+6Aoad8nQXq6S4iVyM+HuWNVq7jwjm
iymF6yHH4bgOt8ZHq0kuAkjQkCbIhxnAjdu6o/Gzb0gbPZuGzE2h4M/O8blIlRyh1rfLSU08WkXj
4+qUWPJvn2lVJFkkZsT9L42Oo1GD/RfDnDj5Gz0iZgP/GcWbx4mqmyJZuolI77K7WYtfKJLFripz
FwFKn4yme2HO0OwUvxUDfZa+qkksXi4OQEbMQBU+jARm5ZQZ4w7MrJGYjEmCMXeaow7kWytOMe5G
z6vGzoKyvNFOHl0mp1hwLE+AtL0mtIrGROWNVYkE69k+ZN0FrvER5fkRGUa2sgiiidZBYvNk9H9g
zDuMn3/7iecTpD0gZMyaoHnaUj+r7NQ490EUZBAeBxxbbqq83+LGufqBmvJ+yKt469/kqtRcYwXF
dvE418hInDlprCqah1zQpIfVe/MR3D7YXHh+LDNXiu/0Ji0mKM+Kehgi0x8F3lMQsvxr1QnaqgeP
yORISSnv5tvlg8zn2QVu+LfIqM4qRu2leH0x4W+ygV+6WULCr9+R+LqU3GnNOyF5+h4bVRcV7mLQ
dwbVZEFjYDHJAKBot4w/snN3i0uk7Ar+E3XLWr3GlesK/FP4naYZKyokiGiuLsFFxvvhgZg8vL94
bk7bsi9xFkbJ/lPrUWA4xo/ZTFxxv3Fxy4kheSb+2mxsvsZjFtsstO/XUH+W8MkiSjhDx22PwO6p
090SPC1KSiqubV5QVRNJHMNNb18H3qz5GEhbg7Bir/B0FmsMXOEX4Wap/1LPfeO4MPC+34vjD31O
PxEQtU/eeX99WOehKgI2b9+0CtHNE/UG1ly18jpHXJncGhWv3bcwCzKvTdDrImSDZPP4Mhc0+Kym
5SIuf9m6n6j+A0jdV+lNeALO4tDAv9YJ2rgrkI3PraBVjet11Z+beyfelHF+47liCYKtKv1/HSEC
wGhppAmEa5YhMO3rWnuRb/56epkg9Z+kI9ApIfNcp7/B4zyQaoN4Wos3uWkZTxyeVVJwJkiWWL9W
8qg51jVgOL2x/mO6zULmHDUILVkFIYBpwaE5R9pF3sBbmDck6oYkY1dCJGXB4Jyi//IpK9WsUdXN
UMor5N3M6wdbba3mojeoywmhkCXjsm8hj05EHx8NCyGsIsdE8VrVLBce2LbQt2pIUHrY9rUUoCMj
504Gmrn96yukfwbR+6v1+pXjwG+iCVJDvj8IxlBWY4ns8//APpMuiz7nwH4d1xId/JJZPJBA/cAP
HsUKxoFRzcMq+bOVdGlK7cnUBF0wMYxuADGx1IA+O265WtRwL46EJKJJwA7To9hw78ciLgoTf5UA
5hoWYSbT614YHhViGDsZ2t22KdR8Z/WWONWXyqDNCcmyxcohKe81Bx9XIkUyS55tpE3xx8rQA1KU
aQlhHbuIzCng7bqHfmB7IpD88fDVu6ty5yVVt6ov+9noayYHTSdATsoC8Lg+zVvrU7pi6sHPkMpV
yIibJpMHjLk1W+HhfTbSx4jiwzQV9YHFvmhcv1FJXYAoZsRMDyI8xYhVleid776jKtifEtl+GWgc
0TT+0YbgfQMFLj522cIWTLCKlYNXm6Pcz6rzABhJWKcb2Gl2frfDsrXOW3HUUFb5ElvM+ltROjK9
Y3sgAU6SWvuHoW7rjnQD2TzxZ0aK+YSHX6NYPDkIGCpYWEQKxul8FXTtZ439wLV6qPh21B8+AsqD
U8zfKwLrdRVStxBH4jtVCDTlCCC7Y5LC6xW7vTFC3GrXTlEjtYcmrGCasmMAZ51ay8Jc22BakZCu
w821HYKajK+iDlfHQjRHt10gDbhFR/2Uyh+G3sjVjezhI3/klTAXzAfWizDEcamkxqZ9q4N06I/U
C+a1NxBFq/4vwwY1CbaRLDvgzyGRdFm52rMLUj3Ou0AqcU0AOBU3Brj8+mzce/6v7iCgED2S09zJ
p4+666zJrOhPoW9YXu8Q+NX3DVNsgFywAJeM6cUmad5I8N1rqDXZxqVIgvep/a5E8gJju8Vz+Gms
ucf9eTlckv8MZRKbRnu4vZ16neIrYd6rYW7qjRNyy3TocXBAnlW8Ji50yAn/q+GTUmuwOSqUNax2
jXfGY22wiKAb6udoj5UetMSVypsDMTyfaN4hdxZfjgxTeTLIJbmDVpaNcZsKeZmfOYTe+fZMINfD
q6D0Z1xGkwvaK6McdEPv4RqTEB7c1/6y3+0EUtf31wcEOiWL5ys5sIC6j9Ba2IGqSywykMu1sWK7
OsBbgnc0bC9VQXp3Q2Om7bEC6AAyPyIFb73OokfB3wvM1ADgsScKxF+6/QT4YnNJ7i4WK7NWa4kQ
bwPId0VlsjR5FLOtsNwwQJpLUEfHZYaQWJC8fHQYXdo7TrzPrnSOIe4yIirO1+hrbIEgQ1Pir024
I7RPR6oZoUXC/9N6SZrLmZADPhV13me/5s7ZBMCueF5vwGEqtV2wBL2ptVKzEpv9rn8gxeEEo+JJ
WtEv7zBrIvOoJtYuI39eEgM1m5eW726eFIjo/CGFlEFMp903J7EyBVktBBi7QOrYpS7Ze1UoJiCT
VloELXFB4pYkoa7KTHtN+34Y0TEZKhzMDk6i6U3qdtsW3gcNiQiyahSliJBn3vlm40OrtZGsGhCA
hOou9VzOdE0gFPTYVLI0QvOD01wbKliqbmdwJ7BIYc4Ivwhd7Y3poE+/vmq06nHRMvDBe8fShiBb
SssEiRK9ARKEJf7a/L5dPbN7Yp3UhlqV9vhPudPpkYLnC3Dw3Mvmws9m8CCq0WxRqQFGKaEh+iNr
0WYEWGihfYHMz+WKXZjdjC0RBZ69fqSzTNENjS1Vmk9lkDtJrhtct9FNhwDgdI8GatMh0wmOQH3v
SrxDM9P+JoKVlj0czuatIhjFK/L35EEMlIbFBQKZQ0LATSJWZDEh/gxmU9eWiU5ZGNZ75DMJNc9G
bPREwSIVZNFsswZZ6ENgz5/wShNw518DrRyJnhJAQEe0hO8vzhr4wEWi2SaA7vQY803Nrt0um4y5
SPjgxFUXanz53uTamIxm/9gAi7GV/zkpBuCsEe0d7Nf2AI07xTisJmgo+cXv05OUA2HSg0moEBft
zbQhzEhv+65OOr/yPXtg/WKkNZMAV91bXEQHtsKDnpKMT9HO75wzzz0LAGSOof5U9RGDqQlamd68
RWICLup7zjMaLys3oI4ViLux1kWBL7vXQjvXrb/BB71uASGGWS61Wi+hiM9NqdgNSxY6UypR/NSk
3YfWDJXjDpxftnRtX0wLMMBktw151bTKjMhDzLcI1kj2HVq5cltUDBeN+3C8CjZxUpxFgmqzz6r3
Jf3z2Qcb4B06GHpTQfX+mDtCkB+UNXoJ1Jz7LFSg/H8l495TApIXfjdcP3LjF9A43/RRJ6ANvQBO
U8vWB+SrvPZOwX93JpGYGQxNgA8fUZ+XZfrHJLqKkaWY+9AX7qGshFokv7j2m84qw3zdoEwiDLiJ
oLGr4xUzfECMxDvQUF9t6jR3csATe/zq4Rkf0JERB2xejyKIrKz5oU9xReou/KKluH9bjMFipZRt
jQ0bH+HkH5n6+n7fR35xnrzxvKAQNueId1e5p5qQKCuwWNIXQXGQsLNpTTINeEftQ3xARNHShRhG
AKwsKc5p8dEx1vtddctL9mtpdE9tXGSAeGA3CgSr+Ig8FqpPvIaOD4XWGvS8PQOcB9ZGtoOiYHG8
Um4i6gRwjLOxgrD5YN1zeQBmVOZXAXdL1J/HBX/cH2ll/NtnN9MClQWBD9sHr1tm+jamkd/gsCZo
2pVvrZ8HBExJmAe7+m4Tyxpp5lbnmc6QB9cl2AJTdnuGUDHs+MxeI0i3c89gEhyK19YFt8iaRp5E
LHuKB8k/s7U6DOqauNIrNQJoZLe8uZ0kVpAjzwxxHK5JKz4/Vbl7jbnv4N8K0UaJkl+tulJy8865
hwy+Kht3221/P4QktLxcbuUrWTbprBc0+F+iO5gbcafyFYsL3+gsY5dweSHa9dDqD43qmpgJUMnf
eNBhdTDr4QJcFP+di0DDXU4Ko5Ao8z+WRtIfI2uIavUoKFsrar2yk0yEPr/lB9Fj7UrL7Geg0ppL
facA7lShB91Y0An5fLNu8kVRa3KfZTvgPrg/5QyrwDzobkcMrhhfq8gjSxVz9NJv/D6lYN9Uqq5q
4wdHUiT+XFVlGgIpoUneOSlpPefvdQbXXM3tD+jCyfJJbTOInHk7RbSdxEGuMrboh3eFjWM1j8Ti
664VPO1OcqaJmkCtJ1fJ0lHaHDxm4XGHNCrhc0ghHWJ+bHmL0tWyT1+jozZ4M5UksdTLGL3hIfEh
1IArnp1sT8sswtAatErprwMSupEcQYigUR8P52S3/zmk2HwH6UNJx8N0vsKD6+quo1TxYAvzEh/8
HXZVzu1MbhmSCu0KjgQ7JFngRBHVPgQzR6s+kkYmHjbV/blvz7kud2mlKhCH8jXu/Bt7BhZs8sUF
14zKzlyGUb6IRdO3Wcua9z7+QEnnp9dBmi2ptg6NhtMNG3rraZWNWYGCOqMphG87z/2dagsx3/rN
IWN/CJ9CUToe6NkMw4eWsus0qVbxpDwQfiw/2qxTOYW5AkUw7HJZgO9d+hgn62zWOb9n83w+9euQ
9nrc0rFMAmP9bKbfaSi6X5TPUCu6nSfMXpySpOh+4KKSUXo2oezKeNaAvyPswYkaTsw3yneYl2aH
Y8Zo/LUOT8O+zbpSHitjyTfIWCv75tdPQhwojog+iNPP9aqznE+Ny3fzLZcNqhZX8joFYpiIKJGd
/ltwDIpMbQE/c1ZWUTgwCB775w7PJLb90fY59j86qfYKO27XizlxTs8ArbItI6tt3ZTdpkOVzkX8
FLeeAmM3r2bVH75gNWk3JV8RIg7VluMDguyxSC4xCoYCVfhg9M2gJPRAF5ibsg+uoYTgnMASljLo
TfD6rzdNzdyHAfu8f3tRRSlebYtb8iffy6ZsdACFy8L65sYq27q0WM0hwdelE5t7P/RmWWZijkwJ
kpHawjPCY1raKLCO0TnB9COYmk/nv6UPIZggQjGOLbljRnNOHsnYtbIC2mOhDgWw29D04o+IUTf/
c22Zy6rKQM9ofp3e36feE91ph4CZdxqt0URmfIeNS+IuJ8qVUFhSbqTvlMlWQVimn8kkwDeQLzzw
9gjCojD15Ch+CzbJu4MPc8Og1CzMBbycdL1+eq636pnJh9Ddbgxyujsck2+IgVypFeI6+x2PJ4Gn
tjpfc4Vf4zvp28M0YmLPWR6smGFte3fvTjXQdknLYIMnxPE9DwLBYQcqZt1NR3xVkNXlPzDSgExO
m9Ile+qu0WKJg8SAztHLDoMNBbZdaSaTmK1yUJWHinDl9LPCNm56J2duD9DKy6x+tuy9KIbw0a6T
mvEob5Y7HUvE/zHUL2QX5eU33E7Cr6tFp5kB5LrjN5KJBJ7VKt9EiJSNAaf+InKZku5urZ6q3kid
xW40RLqh/BD8PkjD0idyptYRD84Fo7BeEGM/cUqtUybjRgtxuzXdn1J7Z5bW2mGlJPe8V5s903PV
v/5pClUXKtVl4IxoAZZhKlW5oTiy2b+F+wJyPAR5zj7yeLAC49Q+W3vPn5P6IFU/JFuYQSdH9q2g
sw//QKkheO7p5Occk3G2ZT91zGq8Dgf5zY18e3fxLtAaTu/0vbs6VrukYOehvuqR4uhW7rLxPiMM
y4VFFzClUx3JWSRGUHN3wTviNFYyBnkDuZBYPpCZ9+DmWCZNvlQA17eiqkmi5y+iAgAE/q60GAgs
//u0uZhP/oG174m1LvQaA1AGeABURfdjw1e8XT7dDUjhcE1Ej6zXAJ4KQMo0BkdIMa2D956TvjeC
tgWM15PsBc7VKJoY+tbNQl+KvAawAvjMyeZuHD53p/38d8O+K6btHG0QWNMrxkQTYXnGodu/ZBUH
lG8lCZNx+LOmNt9WctaK+LvKc6R2NFThqPuL1ePjsWDNW8q/LYV3YbrkFwda071pLmeM5vWnr0pN
f19656aRmOr8PLtqdmgP1+PSTg6PpkMW9zO8O0qCX/lTby2y7vhPseLCtL6eFsUPazs775esNdU2
VxxK4LrVKpLYS+bgXnY8NVg3RbiWn7vmEBgPjD82bAInkGEyhn/CmK4Wa8iF9wzW8DD0Da3kywB5
ZLi8AZxRvNc55cStU7k0i7SLaMvSJ4muretmp6XgoFXKfjdeS4HdbuxQTrQuGt7niMml1T1MLPwt
xXS1TozN5J39ds4nkBnHEjVfVSRqquZrTqxH9gd5Pjmv9BzqZ20i2wx6G0mr4qlUF3BiMFuncajB
mfvcI5tr/2Y28ruyH5qUZgqltp3OwY8Q2TLbyXxWVbRQddSPiezZx/VFEKqkwlhDz+6Jjtsr4iYj
TKnHeSEKvr6vzzRQeKOYONFovcad2TgSSluytPOc/Wcq22JlF0SEJZLegyitBbfahAdxrxl2ZV/2
xhNE3YkFQwL+xPiQWqXMu5bwj8c8K0DCbUbXQaO1SUx0BwHUrx28ryl23d3agxLymbAJtpc1B36S
vupxRgCghe2jeOrtQR6BlWtpmD3mbCzqwow+4If4fOCQk1bl29B32iZERe0LckKS1IuX+zfL6gu6
BBGwCU1FqcVQ6YifkVpyEmq7md5boEwUJxDlu16t+ASLXTzvDFYUkIilKqQ8Alqhr3mFNOcnkDEI
XZgFJE3ZYGvSjd53B87SfVek4XlTVDcHUTkBbIkm0IdudJYRWcS3xfHFRqZuNuWx5slzlnjrtOjE
1v8zdQHc1TohD7Se/QV/7iOm5uFfKsYpEteOtxDj920VmnZhzRHp2uj2/S59jR52uvxi1mFSdVHY
3bqqpVF6CtVzXyvhuIaCKnDnFcX5PEN7zr+KXnT/OF+qhda8m6ITyXPOnh/RcAEZNae3Yrs5OfSN
dHitEzZg9j1A47DYhgZ9lhSK5wVE2s8BsAsOIv6qEy42pgoQzZdKtmZ8g9w0wE/iH5ItEWL2DKWC
m7/L49XANbPzN2RZvJQO+uVtA5l21TG60kmdxw4jrotMMjcVfuf313XWT08fWRhv0+4+an0X/p+C
yEGJ9b2m78yIfPXF9Grh9kVRezEFqZb6Jl8mfhlLEbjihP+pUGAGV1xwp5oOrtmeRevQBOPIAf5O
XUeLQfYmAKvtbj1Ege+X7TtnTmhKwog80fghwAjhkEIUypNCExvRmhW0FeahjVGTd3NcLA/oJViZ
HlF3PumftoazMMVFruiQ/YSE4amUd3KCEXADNYEe/j147C/Kb11SfeesozfgYIcOWuZC2IiAT59L
LI6BbavHmVTGel5YXLB3NFbHs/23qYXe3sy2KVO9Tu/K7zavpAyuKooAq6g6Pwj/bfjomAyxXVgC
HB77zzSw9YG1dL1uGLLdbwcgtWXS7u7vfediRHY+t6Ds5dDuHLxLWrasiq6F7HGXtmdWowVZ7a6g
kISRGx0qrLmJG9lEnbssohqs9OnIk/2+KCqEbSVtPmPFuyQ7DyX3uXBxdds9KmWgSyd/5b+JTKjX
0KlBOBnymdlOjbqPU7dGJ738USbNgrOhi25cQnUfzS6LHaPUYQMfxrTSSMhCeXPu7Oot8Ja/+axO
srh5foOkEGnO9dCov796T+rISAClH2FLrM+ZE5M+/YV7CFqAsRF1sNyIAHUwI5HsQyvAbfaP7jpT
qhZlOX0DODbLZw6+lrBEvsPbb21cYxUKNXLf72ZXJNCTbcDE58xR5s3tm8lK1xgfQGl1r6hgRtHt
ggqcxWv+ebO25hKPRsGk/9NfzVCOcZ142LOyJ42CvZn6k5wUolfGm07ItqHoi1MrLmF9Y/Jzt3Rh
/gey2zuhLDC2kVHyC9QE37Ttq9oU+WtpB5UNF2lreDdsPSieNEKTOn+U49VARCP5hI4wWfeResrd
EutZFWB5DGy0NM6ogl42AoGWzP/SKTNgtoFFEeVrh2Z5skh2gBk8sT+gpP042wNjvp/NgyplX2SV
6yTN+WkToWBxsMSi4JwTPgzB88O8M8j7WH/r5u9nEGwLfsa+y+MtU08RbrMa7z/r0un6AUmTCyu7
6dLRZCmw57H+rWJOkMuwX+wNc6H62YIENnP/xK6efQtpZ6riz9hLZFmJ3s7shwmB+BkaTiFJzTvB
Fna+0B955y7PPm+DV9BjAqR7LjqjMFgyYNZBqlmnGh+CMlB6DRY+AP3naTX1aQzx+2hil745JGlD
4DI49diBEsfcT9E7OjwH7MaRYZbK82vTjSrFPDVZOhDO3XQTBnuD+hNjBMw9VHKlf6i+2E3hgGmF
SYbB/ALmvpYpj5nvPEIaJo+JWgiBuJg0/H0V8B6TGaby0gSnnfL7XDj/oPhE7fkJpRYq9V6uqdMC
Zr8TRCwGU81hN25fTXEmBCQFhHQcGxUIo0UGR+jo0ohLihaejLxks/+ZsVgj9TaQ0XXNwiOszpGA
5HKQGoXvKrlaWle4H7aIa2IB4xEXKHOPU9+8Xp7USwM8tZS7uY5tGlLMSH7eXUPV0CsqiJqmV24o
HQDdl9Xml7/q+BOL0CSKzzMrA+XUD8ijW+m2ff2e+PNQhVysxPlmT5TZ3zAkwUV++0wU5g2MsXGc
oRukBCwdxsBdErcc4CSw/SFMzh/GAA1ZO+Y30G8WPeJKvnZTCvnW8vWQvQpPbruhLC6AHgmEqInl
yUqKrCkw+67CjLUUCRuueBlZMXIsM7tVi4iiPHPWspbOiM0ogwkESwuj9UzkNrvEiPCePwNCW3yt
HD0GZPwlLW+ZriklELTkAAv6g3Q1kUaFOBBG7mXHH3p/8qvrG3pobOIKQ67m99AdEc2PjBlYbbDe
jsyaW5938pzL3Ul1MP68+SArGNpjNbFIxVKI2HFFLj+XEPrB1oW522R7bfZGJMcjiye4oX3+I859
GJHvpGqTIjAGMIAV2/UBXAD/XfThZtcDo4IRj+mrnIgcRSYxmpWwaNjGWpiAgnw1ILbD2VzAPi8W
bCZD+4AlFWz3nm5JjRDo+YFDC0w0AN0mDn3Zfl5TsrLVQwSewlnST5wV00lp7Y2tH9ifpLviec7j
YyI3CRkgro4UOfrDtzKd7ot8Qug1NPputvEodqQpsPk4kX+WUt3IlrcAruMF7ZVhS+4jD7xOg7vv
sL5OqbH08ghSdS3MgKMY6WSa7EsFhdF19cg/OPmC/y+VJCUQzwoGGRksT/0udDdFBOw0uws9hseQ
4V0smlOhNKepiqod9FsVnvyqLhI9i9j3y6Gsircl3txE+4/dDw+1t0mKQqle/e5oCpWyEslxoHWB
YCx71bZ1o8NqMZT9Ama5k2+uQpITc3VQtl84Ji2SrwpJZRCL8Lrcu3pLUsxMdW5Oss1I9JjIDTxE
rjSoQOba4HvmSiJqH9JAnJrXfpDIvss/Etf5lqDFnm5z24APN0QlHqZhThPSo7NhEYmb+ew48lrj
lFSJV6sHMmVslS01lTXoeB0dF/8/XSgug7Cswc7gJ8NfwqEyeuLJccXK3mojd9lo9cLX9NJ0xWq5
p0bGHePfndWtR1QTAfW4x3IYJfsB4cXAc17kelog0YElyKN/vBJ0b4B1C2Rou3JmDvJOW/EYO4yu
hxmm+NfxV3swEsAlPnQ4P5tf5wPWnOJaY/fOiUqowFL+GFG2RJC39FYIw0nk4QildAVkFM+EhFUx
sXSsg5ACJ7C1KL4uMRTx2tqPG3Nk2PN+bdnZcaJIncpg5JbBy6AHzOSmi1saLnj2iY0j5VzKohx6
Kej+r9eIR17sU8VVaYrbqk0uUkGJk8Rxdy5+LZYAXQo76do/DXMnEg3Ad3ear60E2o24IuJwRzFn
FvurEYrN4q4n2vPs2wJ4d3y0/DcCwLSa2/I1f4Ko2uDz4GEUBjUssamXq3+Hy9ZQ9u7+uv3qxiId
CJefoeJmqUOheaWa2k2Xc4qR42lBW1Uhme7VnywZlKpXZYXwARz/2tKGM2hIm2KdsU17TqHuUFXM
a8MG/ncQmCXvPRQltCWOzFZrkPLeGtLlhr0JWhwLz9aI9jEYDg4lcCmtDPWsedShpUovyIKF7hVj
b4/zW+eTeJjK0ACl+Mt5KjoSyko9SELZfx4ePSDCxMv2nSQFIj7+tS1z/rZRjkKOe49Y6xOKOL7K
jE8N2aCWNtQZJNVdKD25WCWxK7oCtuevORoI4GOuvc1VpTIAc6ggVuDwm09VM9QEA9c+ZeX8+N9x
UAK3xSUqB5HI5KRhJNlYHKaYm+SKfmsPaI03k1SW/AV3bY21VPoMWtfq4ijUIHcZpcqlH17U487A
GP7LK50CIbBta/mBzkBGwe0OYdWd77S+Yfn2HA631IlBajG6YonZVt6BJQSuF8b4fH4od66lqDdC
+XlskYrIjSBsmbwijJ4sblKnQL9R37PHi3ysP/P3Z7Uwu5zUYquFrvsqu/vrzue1A0CuXKNncdrd
rAhxFOnqxEWombcL3XpQyZwnws8jFKvhVcBXGl6TcuCnIG1G8tRdfpskDvL6a9KmiMV9cD/Qlie2
n9Jf0rJA7Z2nInmpkqaVLE0PITXLskUoKOVxM8evQSFn751FAMMIMncrH8Chowc7jPfqqxb7V5Yw
lxVGahnXzAF3cInWm/75ExwIlOju6fFGqrzu1ehiyi7aO6CTnP15qWkf3ypRGiElqx1f0wLF4cjo
U1xRmwHwnGTIDjkZG2jpyyXLpnGSZUw/8Cgw1SAESQsiX7ShW3ZPrSVYLtLnOttu+7wK4v8xLzMJ
Sqkj7LW5DZuIS+NOUz/L+DMxJKZRUzmGpWeqIOmJLt3KZsxjJIiMkI95VsdARlGme9czTRGBjxpq
mG4VVUsKPsg+MCGrw9QBPPcFl6tfyPgV6V05zOvoLOTy8In5Od7UDyqC329Li67xks+Z/3jQGXSn
cpNW4c0OoCHR/q5XNBFTjrIRhyXtKLeT/97LpCY95cN42WRzQ9PQMTQfvhkcfcGq+pyj14bpnytr
UH3c2NUWG8NhqJDR47TjWM+Nd0JrP+sa+zPmXpzViy2jW4ZEppLgtvL4LryAyPQ2yGp1ZV5SF32o
rxctexN85pWf6Chn05nnQsuTO9RhEunkP9L2DP09HaEYLoE2q3/tA47mojCEsuY/lRBeGjpb6unT
poQ9AacmoYztyz6NiJ2gbe2TPzGadr5jjIWDOJB44uYt/DmUUU78lxazFMDrZfvfy1pLArWBzvQV
prPmyCrBU4jCZbOn3OIQdXDASSA0caZYh+CdGqn6pl5m9CbnHLctxaLIgXZ1J9zFgkj5yfN0nM1B
aJmakv6wgehCX5nTwXHTAXHLQ8TNUScfzssxxomi5JSwwDBmFDikuMP5O6LadYc7qbEiCzw9hNKe
G4NKHUFMV+tI9tx+0kVZX+nSs0MqBkMAcyiRshWrdnCH+gcQDXYDp+9Gfdl4JWByolFRJVlGUoeH
rCw1n2xdTAJlwOo97K783/MTfz48bbKgtDdKuZoEoxWC3rM7tbi56js9pJ4xVbQdHGWTmaeHHv0x
0jIyV05v5Zg9NpA2uEKm/zWeHT7XvUbPZ6oCkWn/HuzpA49QydH6GC8uTy2kyJX5Rb+cFk7lhy2q
y5GL7gLdg196Df7h5n46U3BY21yFayrQaTeoqDaUvnxe+bB55JG2BDSFVLXIOGLzcgLIw+XPU5LP
edM0+Whaha/7ZC+eaVvgppDNlagyRZKlXiQaDOB+9o3dxV02yrAWLLhTHpIiisl6j2zPp10g3774
JANvI846Gov/e8vc+4E8X1xgdu8DzBD7mKx+CFm9+9kgmV7chLQqYYMYVYRSmugJZc2whsEkKFkR
GaQRTcZNu65YRGoaC0WMm27rZ1TjTJKj+lDFyskDlLW7Vhq9Sad8ippD9IgCD64b1vkUyqluibSj
WmYMQbbb4QXynxJ+yQuPTNEw8uHYLSrSfpb/U7R/sQ1VehnzhWuDs4/9LLBno2uifQQcrOtNiVIB
zX0B3CPbnjjWleHsTxnA8/0lvYiwsAb9BbYJaeMcDKvUJLuAQ1kk2/6zVV3qKxxm17x/NLqzciJA
eBs4FAHow2YU8aGblkRJqKkq++MISexKK1Jyz6Fs4XJoMhsgiCOvxSQsw7KcDaIqylo0kPwEP3/W
F9QANCf7Z366YXlz4g6y7gEPVrsXZwMd5Kse7QGMJal77eotBcTASE+qNzopOg1cdJgKzpMz5hlH
SldiBmWiB8y9y0QE4cmPV6O5exajUL4xMabNBv/wjMXSLAL5di4s3VNJUaNms3yM5FVlqhnPlqM9
EDq0FU5pmyvHUoKXYgKB5/wqeXvrAbkz6R/sES1aCR+Bd9fj95rPbYpADjkEZ4LtNCrcCJ2zQCFp
jEyZ9QOBKaeJl8tGyVJ/z6gKNbl8USbjDFIxuBJzz0PxfqFNqL5M4lgwIiy+f7lcKogT+PnZS1XO
727FOM2ma+SMK1LMCLubkvaUnWSgGuHH5OdkPhQ02AErNx5swlmu9VAcchyaOLeIsnqM2rwUyGT4
0UyqAVFD2LPctzLiBn1O7wqOG0QNtcibRigov2FjTNyyctSJyV0bvNkORVfJNPbZFWlNoRUff+XK
s6ahnefjDhaEpq2LjwwWa4LgNSgjR8lyzn49iTpgRC6RUXYlF54TMszMY6v6kkebHsuuMHYVOcYB
d0DZrjD3xbka8p73RRZybtxOYaxI0a6rVi5BuZelVsgkvnPYIqpuWuoueDUPSMUY/ScuA9xgOwC8
xak7BOq+PadKxnovWoYB8VgSOGr13yYn6332RErLwo3CR0goUO2gtiE8h1kej9HwUuBHSSy8q+PV
KhzOEkQ0n9WLBPCQQ9hBebieJ8JVWgsL+puWC0/iDDLnfLmpc/cr/jr2XoqMuun+XuXAtyUrBLx+
jm2StlfZk4idwBTejCNmJmBxdbFvndaEmfUQQp6ucHQ4iE38bW4Ea3FFhSA8vIqq5KwzkrMZ32wZ
fA4w1uqauHxZeaW76uFWnXEF2OyuXqxQ8LDFEy8lEIeIRgqsxb/2xppjuMp5lXriB/GOifjhxhg5
TAiLSrVDNt6VKycRQKeBTP/Ky8ZE2Pti+Edjj6XA5cGiID5f6luhMsp3aHaB+4Szu/dFguoCRZkb
KPhfRkwiyvX4ATzsKv22tv6YjZ4yf71CAarCaoTmuPkVNzENpW3C3rk0RLbLaglMpxNUAq0NlBwI
zY69/oPC5KbHsOeQreHyef2TbDPcJoJ+/S9NhhzCVkCKA9JxxsUTsEMxPz/+tftV0A91B41zS6t+
Kgqj2wi0q/mHst332cfQ46IbW4jsfhCPn52S0+ijOnrHMGrl0wAxmwyJkVmVNtOjTKn3Wv0D/PKi
d08s9/MS89fu9ObTNfT7P/ST7c3ztMY+zmW3kA1Kk4N7iDS6HGoW/eCbhtMkkGbLV/8cJDsi8mFf
lBnFXPtyYkUTVOuW4ns4QXRAudMX231v7zCmnHKZeJzURtgC4ZqJPze6Yw1K+6NKx24KQTTtNh3I
qoHXidZd9gF09iafOBJKuQSbXwjCXd9b/gvcOmFA370SINiDi4qC96UswDBo2p6HfHhB7tnE6b8Y
35l6KU8USO7v64c1IuimtYQs3KsS0aPhG0a+rkWUiS1xgm9MRsgw2plPe9zeeASycfd3Ku00N8lY
eQ59L80Bq1PTZa0VqDZWHQUNfCUxjqyMZ0xLeyO/pLBkx27bfIMH1SQgHanULHbgGkGOiTyfef6c
R0ra+TrfKUXaCDtn/ofdWrhfppKt/BBj3B9SVWkurODnY8DXmfHUoAMUrmlAi9v46LweRJsAXKIu
2FsAqRrEvwnv8tbRilrqfqn4jzxCqQkYjh3vtJkJXCxxhlZ7KpIy6X3ymOA1OZYixq4UNoBfDTNR
WVyPKv8usUZmNLia8nYhosUZb8IZleEBS4Xl6/9gNJHDL5atBf3gedrrNPKlPinYNevxc0hOX5cj
m5vE6bY9TUditYSWEQfkIYtulrV5h8M393jWXrYFzqd4J8DvtLexg39hAvAD+3/nob7ijDQ+faZE
G3JwQUCJS1kcTiNsQI9p8wuAID5I8/lA3R2fyQn7mER298saAYeu1sul6hpRRvnIEO61di7ZOb2p
0IaMPMp8OQammrBwdBs1lXDTGiY//L1ptZg9NmXtN68tKyq8sJo+DlESaDUrcqQhu3K36f4dslM3
nPjZpZ8nGj0CczcL1vZNcY8fXrs1dUcn5MSrRpOmR0StCgeWuCziza5rNSRKvTtSOZvbzA2rD9h3
AtxyGt3Z0FGV5U+gqtL6g/gSRC0gTuvnnDeOZZbofrj1VkN21miEI+dCqLSynCNx7UqpNhpr7tRe
bi4O9EpQQIt1yLLWRdiIeg8oTJTm9kB8XBoJBgCETYyBQ6cVI1ILoJC0DJJznB6caA4/pXOcJy/i
3/pWbZnqnBCHf7DXu3mig7l9wnoFZeR3RFHCbScogKC7SXlYhCgi3SV0QJcqm9uVjb6FWMYUfXtG
wUEpjmukBHdDHvp5aWTLS6WBoYAmXYAJKRL7MTcAaWOzYqwEXJKpfM/DeGoOV97rsI7466Xfvelh
aSxG1O5z+zLDq1lijoqbGZrwovfnIGJ/YcTZP0Da70j4XqCIXY7XfqPDKwbfBN15y24+87TACWAr
LbRF+VhAYqOM3FILMDEylMLhpRJGb9jbFb69Bpiy5YjxTcsm/FUOzuHRkErDyytkqQXyOBKFxwGh
9nGYAGQlAjbviEkgY/58JQ0CpcbTwPNu5rHRgkZBp47348IeV35+4X7br/fiZBlRZzpO6QnWH3mF
V8ZjCr7kErFgEdaBFo8Q9ahXdLn0Ed0OAXpmnpO8Siowz118uCVNinVRXRjAL+L3+s8N/oKg59qg
pXvLWPAs2gQwqHk+lkskLGwac7raFuKncb8gFvmm2EzAN9SJJ64nJymYdTktdj1jQ77SC2sZqRPA
FTxzGulR7nbuaI6dIsbjVH+VLJbjbm/LfmN2uJZ8734aBRO1faOQR/Fv6dpnVj4PH7jBlc5mcDn2
bFtSCIxifqboJcAQlvlej9OrBkLHYpMyzLpzJxACm4XjNA+08oUIedGg00DMcY7j40ngnDefv8KA
zDEl1KyYC4Xr0Lrpcxa/k66/MoJC3S5DdMbQxsvBnl/g1UV6zZlIeB0PYLbJLMThJNeT1q3mK1n0
XballYpPuAwDjHPZOkb86rWXVoS8FalLOtw0HGWXlfepQUmxxAFFxiXdQznDMV9ikDrT+xKQza/C
UrI/Rd7IocFaTz0KQywGhy6nbTgy5Jklg6Z5ayOVQfMV5zRseGyK1lcuBpZtTgDCaxjS7TGNQh5n
QriynZcI6xowUrx//d53AvzFoUNaxoDKvP5Td3s285Iqp9HXveiJoh+6ToPggYVbl+wa3AROk7QY
hA6i2y2XsRrw7nfJD8TN+DCw8ApKgOcfXJ4iH4Ai+WCOci+4PlA0PolrYTBvQIYaWRwxd2rUdIDO
MvdfGVTDyG0VKEYm40iWcrj+8q5ey+Kt6BaarW67A3VpqZiw0A03WGhrFHvstURMBxpE7aeItIrJ
IBMKGxYYaifbG9bEJvTAsjt0RBGOD/l/0Jcdz3NKZ2X6h7alA4kovn9u4T2AHPto7+dRCKHirPej
LJvyNw5XirityH7mRhqIypNjQlJis5EyD7RhNZojEdA+ssv74pdrARXf3b89jKDMWhGaYTgtPSCc
l0B9RyAY79ZO+eWFSisS0PxQHRCGQawRySqc0dt3gAAzdGyJuKsaiuQMdsmnxTwayUsl8NY4D3jn
qPHd7UJSBY8JWF2cxS63F1ptTKdDdcEpP0X7JKm09P/DR12u2ZlT23slvAss7ZBl5Q/t65lrEnLA
PTPzb4WJhS2IWG1NaaklbISrVBFbM6+MzKxV+eDxgdBV6dIg6UWqYK2WSeSZvwv1Q59veUFkXul3
TJO2ehDeAix65qpouTsqjwMungKypRrwlsAklMhTGK7LR8DUKA5oLrotgLvbCKc+lBSbqtARFx9F
a/4s3akxFFVFdX7aCT43YFuuMxUiJuSJIu1iAJYYF30R3rjCZVBKhvBgtGgp8D6kLkawLJgf5HfX
XYYQ/uW2rkeKsPuhOKuKcEaHjCyGsksnQaI4Uv0uIWqgp/9UXziFoyQ2zPQSYkQ0dq0L4cW1aJFZ
bVKMrVSK0n5a92vmXIhA0GpeANGyi3f+MS0HFyxtmrEsyh3DbdgbhYfyE/0M6ZoeAqUGn2ETNubg
gS+bxCgM36s6u/o2ZnJjSRRquwEhXTqL7mRCDYQ/Y2C8KpKHsQquIFnPfiRRhxfevfGUHPOFjZLR
5ceJ2ST293LUpPLy36ZLeY4SVJWuxB2Yna9ujN0cFAG/x9IlGV8dlWfoJsf7S8fCq5haYGYL67PL
+q+hubdf2/xbPltUr99G6D+Njqvvnh1BENdfhamRoc9oXy8QK2Gmw1Yv6kl9hM36Vv5dyUfyHX6a
CzHuF6AifdMbhXcke7cpzjBDgDOIfvWGjSX7C5/I3KoSBVV3JqwRzcQPus4ofgcIyEi8/lNS/lsm
Fq9U7Fp51SlFy1hS4uDhQjlPB0F6qM7b5UJrtSBS5GXkerQ03WAXK1e98leVzBzQCAaXA+oDbGLD
ynzxSNmaBh2FfPRJKWxHpJV4lraRuoN+EtTnWEgswhGmNnUqf6ctwiMtIVPp4dWc2MjvQ6kZQYct
OjSCFy8/NRi9HaQ36wPjiVBZImJFvhEtAndqzoZGB7CIewWZEea92LmDM1dxCcwZGsR7IXBavan4
vi7AIGITiw9qRCyS9/T8XMzmDcUrYPEHuQFFtUiAz6PUvJrs5l5nqsxxqpY7uXxONfuQ1/zzcT+z
kWaF0szs4BdSYVLyUsdATSdxSZ5x1abnPAZaRQDeAp/bAdsfXNypH1xY4RFmneGQoczsOD/MA2iq
XzJNdo6Ay/SpTq91yXpBk5wPIEZ+fgsuxzTEB1XROqn6bd0m8ZZYmwY/CYPoeDFhHmCHtgwqClqR
PzaDeMNYNVgBKsE552ngGOtMoDpsb+Q91IxeOSW8TSSC9BU3am6fsKP6YGDxF0aUY3nFjidPdz+M
EjOQVskr+wSkePEkOyd9QQIduBcsGP7GMgiS5GRDeZDAan+skxQ3MPtY8ZHtiYU5wc53J15kcXSg
msE8/7JH/lD9o3mpZCT24/4UcGGdlL/Aweyr1nK+4k4Zfvg3vkbyMjbcwDN/gNM68YykLoFoAXjD
ZjssO2jmL7Z4U/Vtc1mzaYDxWN2etW6RqdbK86pxbbuafb6HzYmRmtA0VMa+5kAHsjNmxy+fMazX
xAf9HIxqxavbectyaaCQG8hNHMUHyuyQqf7IyRaCEVADBJV+gNhzNBfaTYN0sndYhQcrriSp5mIM
3qOR35pywoT3YAesb5ypalsmKmSesQYu0RMwx4JnqHtHF50M7OWhmeZ7IOUyQ1nbKXdqQtHLMl4M
RFJz5PaNxQizmYKFwWbcoBeXi8aFtBEmEFFKvqCN1GbuIKRcqhTPUSqngztLkWSlHgf9H7cmO+iS
KxJnEUNEN4rw+fY+tRAZXZvOJY+vaPeXQwjXs0nw3xO6b+6sazAfVKNX9Mm3tWIGyv5OXNz4wFmK
Cr6HvhvOSA8FnGgoMFL52SmWnucZAHKVVuiqGHyCnnkxcWenMQNklsFms9joSmBvEKiWadGhvBmd
tVaPG03jglAMqinsOpskR+ZTRFGZ8jHdGNOgJCjCbN1zRniEckdwypkakA7Z7zLdn1f7KzwamYzN
gDvWNguiVV3uGWt98Exj9RlhFvE2i/TmGip0kdbuy1Mv4okqPd9y4u/1gVKDNNL+ck8MX7T3KONZ
o0nTNPTfEjqiDUCBNa/N1DpUi/OYQbqCU0c3BnRsoGGSFgItYV9jGLx6R83aOmljc/ntMuFl4RPm
gRtYcqjWLJUPmJYamat3ywkQ2JMwSyfDm4I+WQcbbrasczh+rv+YxPzdooStIAlVLm8lb4AJaKCw
c0fsuPybYKhRugZD0P8FfhpWI9YY8EUedaxKIGVvZM6oLYMRTyuSGDEEZca/3GpFajt965zJlpCp
Tm1uIi6AYhBl/RvDuoFKLDlRrBtMm44pXyMNGvbbjb/JX3RfFAuirj4aIIQJon/9gz2uEzKKP7N5
Dxmy+kS+H2/bjZp1XOPJuCLnrNGpaKIhinNrqQhLGA8CPoihgnsKDmPlStqC9U7Fh1y3+EvLt3mq
3rl23gMXjKy+4//4G3fWFoFe+qtT5wL61flKIegvs9dxfxxPuioCJubZauHvHUiGdTKMPVN+gHTL
SkTTHJVJwJXmX9jtGjoNwAgX9ACwPZ5BP6JsJESEXU8xcrPj1b/8N4vFoXIFdb2EgIYitQZtn5iW
9bbkTScucVPYxMCeby93NBG2ITHfSUW3FO9HogUxTt4vR32hBlAQgJ57PhjHbdXqUW9RNTTzj4dT
3omChyHs+NHvnZuTNl4EYEOixGmHv2Cykc72WxsGCK7XmPrIH3yn7mDYjRReoReFx+ct0LcgFPnt
r2aQ2L/89ZDXaffjUHiX80IiQ8GFYiHSQKSMLowBQmUKe/h0UUqmYvXOzzDbs62OA8AzHgn2JxrS
C8hyOpmAmFflQ19/RqDxOJ2OaEenW5jYFMr4r+kP9qM7RZGsi23u5AM1vYxL4E0+aZ3Co0vGh0wU
a+4ejFKk3k61YfZQCbgLnQ2i3CUbaCSx244PjybtmN8UdQCUpAla2IQ/85JORDz728k3TwuRTS5s
dayWdfT6Qu3vM34/vByRo4bLFrNixNCDAXFDE2Ys1M+ExljzsiZidTpXS1HMPQ7n30ysBGef/CZi
PejBsOB5KkxZDRX2EO1S7Ft9ejK7e08fe+bL0N4j/UEbivpUDHf3kKNuoqUz+KH1zjwwBHCVOSsp
HlakqP3dO8XFYjcAfOdkv0bbQlEorbrD5NAKo0FRWlEemefEQwLM1GtdWAnBczPv1eeHXux+SEVK
VEX3AayjzSuBmyW9u1liJIY8rzZZI3v+bxR2g9yXP+w+K2BR8hhXJLeIMbAQFC54wyvgv8//Fafg
v6vX3AkNrFTNb+w25rKY/LiL9tljTK29IOIJb3gcpNLUT/TWPdlyMwlaGm8yTIBbDYISOBxBXvL/
83lWMrC/vewVxfvES1Mofqdum0CUGDJzfebYUyoz3lqND9f5hnxYu87JRQ+a4BJ9X51P5zU67vXk
+v+k92/Y761M4tbuX/pnGF8Qo16taruKfcGefxyojaz2krVyo5sbwZWr0T3/XNGI/eFvNI71Www6
xZCoJkxujn1i58XsecoEsA/SyUfjZeHQLpo5JduEF9LnuR8ZAp/WOMhgzXslSIZUaAv+9dxVhGED
T0nmu8tbw5BmgGnM0676XJS8vq6slhI/j9YHx73+bx6EJzyH+9fpoXayrQUt3i8Jxhwu3O3v3m3R
VIQn46M9R6rNY7Af6WPNJ9uErmT12jUpDZxFiDfPPGSo5/ozvBiMHExHQK979V0ucUnuS9k858dn
U2vAq5heZna0lkBOK4MezqD1RUGOATDArui650UEBg8yov7kQWfdD9oLPoJYPVAwOYKX5pxt1b0a
5kKOhizL8s6soBcLMlPr6M10+Kl0FK77yziZftWZcUW6HjUVHhgdDDUM3wK8XSMhyvstBgicjYwk
ACtuVCyApNit9miOTowa1PsoQLDmnRmgtL/C/GNKxJcqQHL52y5fp4byIrvKrMJhEHcbsukLdyPD
fvJp7aGSwr0mi27mW0mLfV1E9VEK06uoi2OXSpF/VnUZl6v+F/XRQqNGSttOOHUa9Hrujmg+7LJk
xRok1koW7ngmuVNnKEDjHp8eSRN4mMQ+rG9Pg6oYncn9x/Ltrwi6by4XEIuNS4Q/7AlPui+W/WV1
CWzHhdZ3oJQkkwfeyjlL9zL2jY7rQ8VFxPHULlDygW2sqMRJwix/UccHdMlnIsfy4jMLC4V15knz
qp1o7flmS0ryny4LVogKOZKprE/frSA3wRCp24fqr6DIat4k9EhfC/VB9khmmwEdnlwPgKk4FKU9
izaS25htd9Vo1hFBDjLudIxM78CgiKHeAR8V61vR7lyBvfpgJsie23C0a1bRAuePvsM7hHeMm5HG
6wfVSFGTnbR0nC4LhD+mdXsqTPVEBlp0H0rO2dPxbD3CTCAYv6XxJ/4JeNhYP7oC3TFubGyEYXJs
ttWfMlFsDcKwukl3jMUj8dtIKmkz+vWVNpMGfnsQoDFWvX9U/fl/50g3idEDi8H/wcl89QZNACF+
OVKBTiCSKGiqVfbM6vr8ZEIZOXzkWvnwsIhsqy6UCw3qBqa9NFigPSk38OVMBVqRAaG1ZEG+2I5S
R0ZnLu7uKN9B9vEy/Nmhr9L7KfEgc36HAlMEAjdzDmT7btp9EB2aui7iR02BUOVo378B2x6nsGY9
Oy/Cs9n+Vqu2HWPCYbhv+TDOaktfv/SP/5fDs3hTwIHH6eOs6ZpQjALUspujZtOqqJJga+t+uzh6
3M3ZTSdMxyqWAnEUhkgOBc3QGelIlvYthEQqpvSHD/i3KbBLc0H6SUW8WgjzQRaaUREOmo67oVhj
tmmgF6tPPgaVwxnZV0bTKeaUddbllYpVR9UR6OY/O/hXBhzRbRSQVEG3J04jj/aaH1X27ojHxD/u
NnZfZe0FuAOrIHSc/MbMO9baWB/+RXSfhNFbWS8IvvyjQTF0jpTR6CFySHhzyBkK4UXIHN0fy/0G
rh/pZnmy7LY+7nadcmfTU0sZeRUjk8Th7KBjsrrlBNj9AS0fR5gXL7DhXgp0derw2GwNWvP+GaMx
vyjAh+vU/qpK5yVpObR222KGrOWhHha3WFwYLnwgYAIN3HicCqm0knpRy2n/oupUC9iQTzANyPKd
fA4ielmvFar/26zapABXT+sLDGKb53sWoUkPPRFgX6OtIqq9AqzJZxf0L22Rt7yk6NltjrfDcdoY
sLF9/jU+RxBJvPbhUcNLxOD/3HBjcw6U+GCyV4BJdUWXBj+KYEOjyrtVVlLXq+bhRKcSkTwb2Guj
hWIM9fkzDsJfdvJOwUKLY3VPFWyfUlP4WKquNnVbd4T8D6g2FXmseT5PO5kEmPQzCrwBPMOmWtz5
Q6atoPORGXZSzgvC07Y7g8zhImO1Xu8t0lEu3itB/NpHVEpatgo976t1L93T1m3CN6ovXoDdMOLU
4A12yBD8nOgA460hZHQp8REaZJEA7lrSDkbgpY9+HCnP/KCE1+871xwnsmOkAAa1CYqaQkt/AQ0L
LN3d64Khm0DGhKWMZjpXRm/HkpJBjNRHPMGdSnQfkxNoDUE2O2IVyHyV4cCfVweraYQAL/zpmzrM
LtPKIFuuGyz/lgZKiqylRK9MLj2nbVY/pKjDDC7IYeFeP4LUc/KkVx6VDldTRofrzdIoFYA3+5Ao
gikXpCJw2zl+lcL6F6GcGeK50zp+5pIaGYEJzXY2RS8rekagUyhYDrcA/I7lyIDzLAVD7E4864/k
ACYDcdodEAmjnK7t39hjTtAZDT6ItdgHjT9S6ncFpHWSmBs1RDtTFcs3KOr2WnYN2MV5tVvTt1hh
Qv8BQC0i9OQS2qPjQ3dlERd4eSuldhTr+HcLwm3eU0y5ODBS8RAW1mlYJLGez+mlHAvPh6OKeQsz
C9AthDRks+etp4U57vmxAhETmlshKTXc/TRo9oeH07+f7r4eNu3RJxJUvKjoaIjfP2mxWCAuJzv7
u0Jf1l+lFEKGSpfFhIGL7xATGZn/BP9W3WYk5mgV6wrZErG02aOWEi5CzMtd/nPgg1ANuyHkcqDR
C3D0RYwrvOSCDsK8ki9bO0pWA3Fb5/o1ieZ9Os3I0BlQ2c4maiCuQJwA1d6JqSR2Xdo0jTONRF/U
KBAEeYGhcogHDMyHjlcIRWAx3rZGr07P+CQ64vOOqCp55zEAX3gilPr5SsG46kjr8WNl1DhY5tQI
H4vFfAUI/Lk95wQfsPgwRna/zmy2DijsP0+Ove3N7+N+Gz6GovR1W6QBgsvgLZsmyE29T7AY4QUP
wEoTHO2+pRULqQ2TI3w+MXAUXgD3Az1K1Xl48hufSrwVIRxL8uEWzko+bxylhRJlx+kH6u1RKePa
FLGrr1fjxh5beaLGdj6a+oFLhziE9dr9+Ezz/F+hJnJ8/M11oyUCOYTy1YrCEMvNmPiG+T2anKf9
zW2xu8aiX/RLudHGtFU3T56SQqWLa6FoItfAPRspN5cgAHtIZd9ISRPLeq8SpxsXDK8mmb4sprt1
dwfU4wthGog9pTEaV/cHhffvW1RWY0a57L5doBfOOBEyEEm901Cob0q2BsA2R/qpQEkZntXKBEe4
XZz9BOi1aS6I+komktwW3xmSjSm3gtZ0xMRstB287BxjycMj63McIahFTHR346lBXSGjXprWUhd/
gNcNYBnXhIIHjpCkEpciVIDC4vQfWQp/oQNLnrqCLLa1ZC4E/f0U39P8pi6YFTJCwHb+41HA6OgE
VJRz62vDaIrTeQjAPokW0U/IYmzRrzl2K1RjkGQXEqLMeLfJBBZkaRJy0T3qCgHlnZIOyl3eRSTg
6VovjdBKgVP4b3YwZCh4pXwmxxpy9lH9Sxt8KmjrVXE3aJACfXocAxMWSj+0b4FCw39/VsQCgfEi
N2DBhzIfgZxFh0nGGaDVBe5Qnk/gTb8VpgIwNkrc4FfFXAYIbC9cPRNYpkQfICn9LhWPWXiyz4Zl
yULHZbgJ8sRH7id3RPWdKDUpdY3L2ikUzRB8e4P/zj3L7AeyG6AgPNp9oYf99E8j2zFJsyjbYhpx
1hZBD1nHno0Jo4bOZTVfuki/o3WnPJtCv9cEU1SI1E34VlmrPVQZJS/faMRiAPP3xcFchDqrshUM
iiTlcryJs/JTyjmrqqyBQcTDgraPtHvgfDM7CdsR0IoXRoWeqjYc/YLyMFpMbQvLZMwLfqkpf7nM
VWCoQpWKusJDBlSnMPajKHsACJw516FL7RahW+Vn1OQ6p78ApE/9iWeeizJTE616gu4wIYds9RzJ
eQdljW2WpLcpWcBF206S331um6tHA+tgUhBOPCCZURh/EPeD4Mo7XP6ZlM78D0mn2BE7aHcKUTAl
7dJ3M4SkVMo0jKm2bjnJl2zNga74rpr2gMGvMM/smCNWFADD76Bpo3RRZFexdeRUvaRAjhHD94wg
VvDugsUAMEMzcFnvUNDOjCZKlxuMlyBnUczNJm5iSTHGb+Ki9YW1b24OcZBcqw/+JtfKiIPAnmR9
7gZwHgUZzlTF63P3ZB6yGNNmr1cEs06Pu3n3Ooj1L6RYqWYElbHvP3WmwiNwzFv0ILqh3N4YGZJN
AMpT0WXfyGd9KHT1lwRT+3PcfPI6SdJFGy3q0X3KWDkYJBi4E/P/rcGPryADMSIU9Usbo5L+bUti
q+QzJcrFqq62NHP7Wh2sj+otWe5IS3DYe/WE6hmN3SCb1EtCM8ZAQKl0bex+u0yDyb87cFAEQGY2
zhIR6i1vWFQ+Z2hi8iBEiRoO9QPHaXzfoDrtPxeat6jdzuTQVZs3L2J2pMNGPwSGiAKIMFfqNXRj
Ub50/U6bcbYDWBhNCPnt3o8k+tSVFTaJIpfoaYJ+MGJpX6BV4hnzamhq+vjAuSSivUYG1tgjKFd0
eteFpoBHUtKGS5HHJ1mkXFg1q2S4u4RuAhc7yky89BmIFKoTc6DjQHhhsDjMlgYWxRli/Xr4RFQD
2Jad5xdLj727xRFCshLjTmnQF1+2QbEHA+GTywZAXyPqyd0NezVkSYoI0a0Ea+xqUDMJvTQO26M6
KirJsTg3zlWA/XZm2OPTs7mIM5DDCvmyXFEdrPSq0wERJ1KSGktoGcWVJ04Q437brJXxpai3lZU5
eEpQNj3tiEtXE2nFFHOJ3Kzrjf1nEtoBua3rOHggYwCg7+ImSW4r1oJPNrMi8rR7uFHxcW5uYn3r
MD2hHCuWiI9lj8BYjHrluW6NI7Skzf10E5H0ziNPQ0hdKz9iAVd+4UX26BRitWoL2rCviRJnXoQE
B+RMAOS0JjTs/gNa3YqVOP0C4zXcTphEVNZDyhUtKwwPYBV7Yr7bJ7b2LgalY4XxPBE4FLagMgJl
owRAT8ufcwtskYf8AFG9GrLJ+pKzk4xAnYTF8HGsEL9PMUBsLKLWn7QphehNeih336DsoGu2Zjfo
vfoXDti8Ws64a55UNWMxCg+B9U0gnu3UJnFRRYV+LzZwKXsV9QjfLNyGoc6m6lDeDF4ZKtUfNGyt
7QFF2GlKi6kPkH8qa3t3sPVdQwTdKFNU8Mfck6tKasgNBiSuitwzy+l/CkTMpcNaFGsZilB5PfSY
w9pyzViqHpMpvB4KWrUuLIbeDYf4LiRa9+3zm3HU8L/2qwFvfn2gK2GByv4N7HJINw63e9FJW0ck
cgcv3CyQOJ9+6em5DyfbbjlM9cggXm+zza45IProoPIal4w4tkhB2r2vfAj90ATbx1+Koe6Hbw5U
/yEBThGuDNlR2JzV/MCZq7GOjgijZH7tsBxLOgFhIRdRoSI6ZC3LmSkvI0WTMr3MiF5K91vxi3vf
+k1FXp6fIUN98X7gbIvyMX3H6WLBgw3aOWew+nNClvkRAFHuJkVdmyNFYQRW5DLo1WbL4PXIlRks
dfxpGWOkyBDDld17mRB/WCoD58932knjjHpKwmm5YUiAeuqe0Z7EpmieyRqRtcSKjU6K1NcnGBMD
ir7KRgn9julV0x27cPQuIYKsc0SN7c0MzcWXmvppJOk0kh2Qgjieyv3S6ZFBANZglEBG2LuUC6Ji
TN0Uis3/Qy03graWbIHTPmSN41J3c5QZWAHJChYmklsUsA8JLRRuEGFWtTTaRbxduB+gem7j+jVM
DRaDmtC4eamSj3yuA+DtWrrOuHzd1BXnte1Bgc72gKyfj/3o8+xJo1x9LYCtT8t/8JybtnB83v2d
9IJKY/LKyY2sWtwMhld76udRQLhahex2d2IdTNtWEm/kmMCVXcAh9rcFmkWLC2y63Paqt+uZIZlz
ku9/MLK+VOL+NNDlhu1TNrHS0myl9vYqVyrr6zL3O36RaPunMO4azMjDOc1hqTv1VtDHyHHI2h3+
GFRxMJqqps4f8a86DUxlX4a5FEhrD4SUgy6zkqXOdwZj6ow0MgDxzUQ2zUS7YGCyP1AdTEPcWR3+
eStW4oNDd5J6P4JoYT2IvLhcr6yFrZT1GDWwgqyJGlPtb903hr0LAPqi4kSC6zjxtweRoGjIFfqS
KHnuaub2MnSYZEyFP0VcJEF1GesvSCRw5xinYR5l4hiWhYY3seWT/tT+xq/DQS9d5ezzWpp0thy9
uTMsDMxABbpkXI2wf2SQa0HEchiT/hDBk0NefICf3cQtLrgkZA+7rgmonVrB41a/+mPPMEDBi63U
KS9iH9pJ2xYlwvGVk56XBl7SXPaUfed2NTfQMN/30XS64AIPrJsi6ArMF8ABnwMQSqhJSNCtgrpw
21O4XnJLNZmpYYWR+qG1E9A86rfO96623Y+OoGO7TxJg4EphoRVBlUy2PVLro8el294O/c5VHVA5
4sLMYU9/eTK//AIAkOEe718qH6+VffhSDOlBZqbXi0/FS2/ZkuERrN/tYVSFl87fAOjB/bQZt5jT
lfVBt8aj3OLfaBnXiZUMG6oxBDVNxOEsVaKU4ufGah0aEFQ0uI/i6m3MbJL8qVqhDb/l1omDCZJk
1bZe436MDSOd2/dtzMQla2np9vVh1n//qm4zWi5rkm9lLV5B3OhXPLxkO6u0A+YloLN1qcczcvxb
grBjvhRj5F2lQOFYbtEj4mMJaxIhhvfMpE6Ep3yE+hpn90FOwjp2aDBuyDDonjqe37nySxqK88CN
YJyKGCuDkBKYiK+mlL53N+epmQ1HnH3+BsO9sldDb8GTT3dP5MzGNmt+Pdb3bwDQttN3Kt8j113C
eMdRyy1y3P3hXktVe8lhqW9Jl6dwoer0kqnOkp92eZO3xyHjIlYEYOZtUuTRIWuwusdE26Ph8bJG
oUcCNzDNepIab0sJLU6H8Kd1zluxnqGwmj15SFFGBkhIpyGl81cwd1w+ediszfmLVTzWAEd4gDUc
Vz0itLU/me3DY83nD9Evvun1IHl/CHHQq/t+XgRNEnxaZ110otdEHb4NXn5G5TvaYFXHh0iIYHxy
wnw8qctNW0Jp9qMd6xYdGvpWE39IOWn65OQnLyTmCBXJfK2aUXdN+maNh9lXLZ8g9pUuMGIAHOoi
phRtUkcnP0l5BNlTFwZYD7/2vL7z9qZajcGuhMhueD5bH/hl+/MNWKlxT9dZdOsy3/JgmopDLnHx
8MYV0B3XzKtP1HvZGsNm8XmLm4S1VeNvCV1RnUr9kXhg+snRz+AQ/fTBNE5Bo4tfcYp+947drZ1f
41jYrUx3wMcD9URMokaD7338MjdUceuFpd2Fuh/GLwcYePhEQ7OK1dDgSn5X2DtflkBAbPK69eFV
JMxUhQO+483Mr6x4P9Cn6gzNl9W8Wd3vYKHyfAWibycdpQUHMZjVf3NniKhL5Cbfv/zgaL47qOZN
yoxtVy8zsT5dGru6hs9NmJyH4RGbrNOd5xCrhAsfq9PsRwzGKZ8OF5uOrpmyS9jx42h38xvHKeBz
VrxU0s4L08mY8cEeSiXV1qkmtoSH8P5Yo1PGoVxOvv+lC40wtn6lJmWfBFujKH1VKCY1VplCdBD4
7S19lI0i1cumxMURhg2SGUsOzSQyoXarBFwt9MSF8y6hRR2kCr1YrkKH/qSRIGiThzDnN+KNaI2N
eb0utZuy6KDli6K+A4dFrgjsq/0+Sl+L+ExhEqQEgo5eAxeVnXQfXiAJ9+QTVGgloGbYXld0+NRJ
JzGdQRKUBPTn64+cUiSCNJxNEBW1nMAusc5EKmvR9fQuqAt2W4TgF5Xtp6DTlh66n8MWGkNywfn9
dM/Hj/VW9U750iqKNk694OhTwEMZN6myBkpLlkntLzrpe9grux+YBayrGDfxgI6txGBfd6dV13uq
vuDp7IMdz35Tj1IlhLy6r2RICZe1lsc/8XzdmFN5jNolC8HXWN6geHX4hlcT3ZO6FesDPOENeV65
DWAH8ICGV6pN+sAV63/1hWNsSoLA+UWvPGEhpYGsGITD9E6bmHJFcX0fh42OqKNuJ2u0+Dlg4LeB
VLNQ7DknOWYUZ646sKqBW/0Eo8zkjOaZLYSXGBpEZVMe4UWKoQ5f2ToOVO+7fehtag2qmFUXKuxL
wkeBDL9dk8z4N7qcocJdBsv80Lt6d21W9YaHaM2NO3+b5tkChIRR5AyL/MQ6tHiUCWw0ZC0sZEgx
WLoZtiU2qLyFJQScyNGbYg36yqbDIPYZizXSHn5m1sr0bxLJSE2+Yvj/tidDZCJ+Axy5Lsm91IHD
7/W6nUqo7Jsgw/3YiAupbrYVI9AuNcaRlvBPjEqn5p9ZFoGPXui1nDABxfW/FlFUejmr4J/pvtfT
mXRgwp0GAd8ORAHpfZY1CgIdl7Zt6lTxfuR7iNT9gBGjPmCvAZMj6cBhmJHPDZHrN+SbFpmoNzix
sr5eUy2HoamlXUgXMM/7vlaYKmq6t1skWZlpg4unZZZvqqZp2c85hXLAyH4uL0dPsidyrcUwtX6X
jpxRGNSSurRddxdEnQq91+KR4R6oMFEAkHvtgIhfXMWXUDwLZfOAQiNlFOE4DRD/xqCBIQBQEizF
Oj5VusOX9ZjEdFbrgNoInniH8OaGWxC+hByO8Pwd4A6hZWNsrw+piIj6m2zj/Xm5b7NGvnx4OJve
7i68ERbxzTd7uWDy5VKZozNwiDZLhmAQETkxB7QMhwNE7NRkQByalsAncMQFD4LCZYqTD5Z/9CDK
4sNQYQNhP903wVq58w4E/+gjONWkhvkyCCCtNMkuDNkQTskgbLbtgKiiwWLq53Ks+UbC2lSfLVWF
vkM84P8R1q0uTwwy0vFFlu9Xr/KVYJ53mndG3hyB+MGWuArvB0Ny+47RzWs/CIxX99Cq9CcJaSgY
lroWrjuwfrJX7/NM
`pragma protect end_protected
