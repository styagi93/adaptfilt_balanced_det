// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kCn+ZfaA3MvMq+gs2Dwhe0gtpypTsqxJEj46kDGKmYEs7j8/p+ddz1l08LfunZRh4B/kSCk2xIYM
b9ugeDzhACdX3YuUL7MjXPDIfRTsZOKzSGlFZPyMi3rzwzNEaMlwmjtTW8sm4aSmwE41GBZgRV9M
8FfxNM7WUOdB+fIW8HKr8Xrko/jGYAKkYvBPOlrcIMZnOJAkI2gURVW6Gn3mZRs9jps1txJDKsmj
y1OKrVj9xk6IFaLYzNm65RYGdNDy6jjnhIyBJquCwlK6iOPi3qduucimzC7PdmN4xRUROyIBgdp9
a49kLXrxLam2t3uCJv3EV72USFP8wUd7Ti24Aw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22832)
a1nUoomPeDPS8Cql415lKzJ8BtrLIVCByAT4FQso2/HIJlWReP+UdVjYqG4oCEO6zaSfGr4EOHs5
exxmw8UjUDfpaXnZc3p7tapfoa6o2/mxEs6GvkiSyJGRkBrP+LhwiYLnzg8VuhJkQMLCpS8w5THz
figsUV3SVJe5D/Uowqk/NlIoscyplc5ohOfGobOgxY+K8B411/3R3R1Oxh7XB+dmhCOFQOSerpOI
vSuDebqB1/g9RuSbh3/DKFM0GVA67BFfIDr1ibNnYF9NqG+codulSMWXkAjv3w1x1P6sFg8f9/GB
+mZN3GzOfyGzoVTzZzZBuuElPbaiTtzb7RTMnIphLFWmWOa0WdHebFMQ2lTVal9g2rtccPuxJcWz
X0JyDQdDib7nVFh+AWv6yyEvH7brVgcbBjRishsraOBBE4ABdBR92wRdXjo43FaNEUVIWgn6ylS6
NDe7TFkJmWRlIirLmew9yGNHaPG9dpriXhTTRUa6h/3GxINR0bzApiABjcLfVQE2PRKIFYgvF2Ww
I6XckW3WpAEPhh3Ob1j7lHNu5wlXP9ohXfrpXVjanGQnxwvCAMUxnNrEiI74FeHYc04uT8ez2NaD
QSyTUvDruJAuxQHtTEOY1/V9WEB/tcgUhTDZk5dL5SYcX22abgSFSKbWL86L5Fk4HQClXarC2YKD
p+SAXeSDViYotWQWPAmW92tlTUroqoT05Is0t0oROXZikzOO5ye6eFNElO6hHZ9N262C5aXYmFUR
yerYH4Nfq0GWS8kZoiLeHiyH6jxRcXMOyWUl767JNTVYBnk0LusgsibwbVxz2sc3sX26RAX/jMTY
gxvRDp3jqIQcrtg+BhZAUNiW9HZR+Qv7gkP1Gri9X+QObEG16Lj3JzgJ3pxIQu2YocS0YSOqxZp4
8GJ4+xdPRe6SkBrYlmV+S65yIRFZiDxqPcnKGN8xwmhROKjO3N1Pok6qQgy5Zp4GahBF+MH7sWLw
3nLXW6c59UGjPok3jNfpzSLX+G3TuncGM4gFsCTbtmg67ic7KiBGYyFsDIm0sbtu06yHfWDYQkVt
aaGy20gsWhrA10cPSc8y1ivgmfjN+ftgMdWQlAu4yXs+e9ykZt2lKmmRmRnEihUdlEBNSaoTDV3z
oBLXB+eyEGKxDItRkttl8fdM+YZKdriB3bHDNYxiheHR0NW/DpMvfE+9oHpgHNsCawQrdHyOWuDE
xH/jUUoy90ygP4bybXKTg3IA5gprdEXb20wxDOCnGloBs7zk9tuvD1o/7kaR7ur3gr6O40ZVfntY
yXqY7MBapy7sVdcP2GAFkUK7MTqiNCG6k3G3YafE79IOsW/wAXUL0v/dhiALat3XjiVZjTqo/nxc
t74RR3VYlvOURsnHsg7TsNiMWfeIWlUo1PTKyV2raZikoPzvswWsTSrGbeirV0bxqRNPeh7VUl9w
9/QUhCnGkZ9D944tW07qwROn+pO4GhbR3Bs1cTnwovPtyeFT9/WvZH7/RpI3kPBt/aRDC0OHZmYe
z/fZRKbIfoHMB5dMF1N4lCV9UO6gmgYZD4PNZyAVBaFXadbVq1nuhuDT984dig2hNg087SfjV7Q6
d5MwDxaxFbosEGkSutfg5gVR5dKRYld/SRTqf36h+T1ufH+wq0YMOO7WRxG4xRnn2totgt/xX1or
d4YkSHfD1rmQWT57l3G9228IAWXX4+U+0Ui3McTrY33kHxVy2jDLeESJIpuqbmDppRuhITXzfmUv
2ih+xuZ6ls/diTORf4IerFnbcb4qh30g19sOvAkpIJQGmvwO5uJJXiBJ/UIx3BfQkMdPOggWw0ID
2HJviAFFcUtHpXwEZA+MHKpYKAmNAPuvBdvNiG1W2Ibcb3lRqHlv1ZL6feSv0w6YojNZ/SuEJkaq
NDC3CBfYNRIB2txeQTQFEzO76iCp84Rz5tVkRFWriYAJi/fgdtQth5ZYnUZ7gNepS1OvimG0EnbR
+CW73wFHBr9gxnNWrG+EhcVfZ8MDxo1HZrLY9wGxYucw04siRqKsfj71xCwQYsYR25L5EZuItBAg
TF5RERvI9Bsx0X90sQsqIkaGAiQvf5cpvcYlCw/ltdPV9Zok15/Boga4YCOQlvR9UWtcgzWwTI9u
dxR32jdU3uHH856RbHFYzDc56APCB8pFH1u1jjz5sDugAl6lSshrDwb6rYY3PRMp1eQvk/46rpMZ
nHr4hrwbtSrDuGoq7aCe6w15lGb1rNAkYIo5WwHFiCWWaqqR/qNGRb2Zxz6Ax3M0xBnTVaYEekUs
zj209/sqTIUFqc2eWX7QLZVCc7xOXHYSMzt6lHZ8i8stKpTGJcHBYx1PXa7XjUfQ6UneDiyJfAIo
R6wqEWJhMvoAVc8IuQVUIKokrBXay23CTMGzcM5QEtUwYY1vDFsG1NLxuI4vUGukuYwyPvHKtQ3T
cnT+z9Fb6ub/qIf1f340GXkGaL7dc0mY+GWuM5vi1eiQOqapkbXsOwfiZcQQAKhPw6m+U95RABi6
i9S7P/9dAaZb9XCBTmtPHn0HhivozweYekfOsw0T+kJkc3LDqq6evOx2AEV/6cMlyJtkNxSFxwgA
xYTgbiQa9yK+QjPVXCoFlRPs5TDygKo4E564DmFLORuDdFVdEajZgUY/Oi3DpNENbko2FWB73jFF
mf0ViOqzrh57vrxigmpoYxUlz6eKBHLs9ai9EOK1dyA9jT2+XPsp1fULi4O6dTDE6VJxc8XzJ0GV
L6DeaegPieOGAQX3yCIrpB0ePa/4JcnhjQnFzMXfwp2qm2QoGHGeM4x+ys6i4Jol9PqhhfyCe3bI
mE3FFlDFeEQLPpRgY/cYRr2IivwLUi4RqJV9y79L4KlOpgH65Ej/c77eix7UMsRCRenhXHvfBg17
dq1YguvAwQShBhbDzwfvMKlSHi4EMD1nJZY4S6/bz1VqXyTznYZVkn9u0RiNxnpmqM9bK4P1uaSq
jo2P1uBzfpDCOvTfta9JKj9fdoCwrvQ/q15yUiVISPzc6ovvqbX3+SxKF58ZfJWoIxXpyFjw12pI
j4jBHKoxxORHTmOm/32rJ5BqXLNxZ/hdLSyzReSfLF+nXshz9Mv1jXYRr40XF0zgn15FIWQYLkM1
zUlizm+0qQUa0g6VOFDgJ2ufvRIsjNSnY53uxutKqjDMNuS7jIqdW40/p2aQFUiQRVIIxM5mo/N/
evrBnkf3HOf4G+jIzM+i6vv3bMiKUDxWXrxSdupnTf0YxHM2njMNKTJCevvfSVL1TsghZdnbFxnB
VRS8pvJ38GKLwtAfbLTZ//Psk7EGvZO7EPCKz/QuzKfEQh9dxOfzwGtyLgL0KD75ljZyRGBwVb4Z
5JvDLEPaxWjoNrrs2TcSmDB+4qCxVRg1kkME/3XyEnPXPW2zkIUQbwV4coFduQhxTT5he8KtI5eg
0MQ/nbCciro8l8iFTOOhuJOhgeb+gwAzwt/nFLwSzxpoKDNVpicengjqfIynM7jS50R7Byo65hd3
a3i1VasPw3NdLeBFzGnw+j9C9XJqTeeweHyaNQzESOCNSSBUjzn3N9ZhTxJ3uOj2m5iAAsJWwwpS
3XNweIAwAu2sh0KZf1/jbf48d19p8M0lZR9owAgAkV08jnl8h1rX1/D+AC9jYErfKVBQXKF+2rpg
s/azbbNcxK/Zm5LTKJpgGROuHaRkIYrKxeQn6KtHUgS6WAUnAjKIKUDiEVNgQ9BgZyMV0EVTeg2W
nhIRpaivWysGTAs8sBj99wSW2NaRPeDKf48larYMulIgS1oVgcPA//z8Ubd+qUGJRHMoqSa9CTDv
2bSFHJKGBuH0qSGu1Pb9fHICtrrhdoQdC1KqS5LJ4V472gKGZQ0Qo1Cj5mRLF3SKqKCNfv0X91ya
k9Ktef7lYbDB6afp/Mzfn1Y5rsVQlCcgD1b3xTqpDoK8c8voNcLZrqf9zu1fyxxVIz1y8Xt46sRm
OzYrK6LEGk9cqYzRPGriK2azeqOj5lweB5ah5jKPDeaRn6rHoUE0o6VKZiUKD4atuRZhSjmt8ZLa
1b0mzoF6bSD/N0n4i3q7yYYHCULRdQA1MZL3CPEwGi8mZFFq9lGwSKfEcPBigjsroM5DlCfqvnNu
SYsZcZxsF94/Xt4Bhh8J6OaYS2eBNvrmMbXphRDxqmisLARIEaoGOvUwHndXaYHXnzM7VEJYSbPm
pA805HsJHXLDQZ9f5hFui4RUXvZugr0f/2YhLUxgqyTWu8C/PLTbbPC+qpXzqu4kJt5a2B4u/gHq
w3IG0FhTjYocJLUsx28imSGoWdZ5RR32DiIDae6ZX+ZO7VkPD1LyKAa03norHZGyybRpjoviGEiS
dEYMvDZ2Mj9HVt/nHi+oS6fIbWs67cxlAjpT9MGug2ZkKCfht0AcS5iP9tYVLymwtt4Mca5D3W6I
CiSZid+91g99JDrlvJLnKkvlfcfP+op3ljftSk4rZUg4OrplQTpHr2fk5JHqJJWeBptMFI6x0kN/
iLjb24zNIYFXG6ETsQ1HG8BNGE8S5Ox2AmhMtGhAWaSCtQRBXnPwfCbpwYEzWTr9C+ck3nVqo+6W
Cxr2QC0+JYJjRQaTw0e/fBB0LUr0XZPf5qFl55q9Dfo4rYIkCGmT04CgCbd0M77TOZxEeABNYT/a
RHRvcBHv0gWBCe0mhpIOeIRLC1oSnlF4UySxnhCJJE4QxKfFrV4PAbUkLNy/wF+5vLPd7lt/D4le
TkDZbtA8cnQPoZ9JlYpNGgyVGZv2Tp715oQt09Hwvkjm6yBecByxcJxv1JqufBO73IxEt4ZlTE49
pvZ6Hz54jNOqqisYsUSq7O4TwG9+Qnh1Kto1swKM/blcQOxOuGT4xMPCx1wFENjvsFI0IY6andQJ
lj/zbG9EGveBNgho3910KC8Z+Peow4vszHi50IUoVNFUWrFqjBZWUBHVINJtbHYfy61jCdF8W5ze
h1RZPBMJsZrkJbjg7gb9rG8Aox7rog5M0d7BYSlmHbstdzgc2Y/7ZONZi0lDIwPFxRH4SuJl+Xwg
VjZcj+QeMoVcSg1CYTd7+4GlgEPYwrplZ5Q94JFWuvGpk+m7E1O/MDXoMzI/zBSSkzwgyPia3j0z
GOkOYdo0LrxBU6IqZMF9Jfpi376tLGJ7P+EyGu8Tsf8NhPTU57GaDqmB4AbHup5kH7U7oXC2HdxY
b6kBDq0vmQUJ7G/Z9k3fZvW2+u1/K8wcecD58m1k2G4xWMOq8UJr8p9iStm/pQNnluBNJ6yHLRC+
RaVgEj8SNlBI+fBxefllqETNzDEDlMBpTBPqdAzFFKWelMvrZoviTyJvDX6oo3hbh2DvIcI/QZ+B
Bdbtb3qLX9R2+bnBq4w7z8Og/oYB+hphT5h7Chz540PVyzRUVONaT05q+bg+uJHvdgbr78hrgxir
0yhcI7bNB9v1VwNzul8eSnyikIp8Ycd69xYF7NlOyBMJiLikKJWQcx0euzgLC0KX5hS7iy25uf+3
48l2iKq2l5SeaQvH9xl40UmMMUF9m6ttq4WhXwD3+0aFqe/u2Q9Ri5wf5E0pbulegjtcMH4V/IZj
fJGbZJQ/95i/2iPFo/waJCKtqcOyTHf0qVUHgzd/Zc+ZmsCF7hT3hAy8CUS0+zlIjvl+sk+zqyAf
EyiO8SfQ+hZPBFBJnq01AsPbOgXQkIx+n5XCs7kSD1e+hUfnHZr9gfUd5FUjd9f1lCn3QGAR9KsR
c+Fo8NPj4PalxUk4vDnR7mfmoDHyviYqHQQwNOL0g4RNR6A1VU5rKQaDB5qCXputvRsoFR9Yu87o
BGm/BLalkYg/YOqkuN6EHr+zsRDQfRyVzIXZ1q1n5GR9xshwnlV4Zu+L9drC3KLyDca9PCUwaysj
H0sQf8s/rxRkSU4Auw4Je/0uqT2Pfv2HE4tVV5HMh1HhEg671m8Zyv6O0SBZXmIOcYPHgToWnZ0X
ljiSDvjD64Lf63NoegI9eYIJECrXuKbzyfz7YrV4NnkzkiDztK6cQ1AS6VBjSeqP1THvpZlcPVmj
FD10319DjRNB3fn4p/oGYzST0NuiN4KzM5sDSiDf+u0ETs9+lPwUalodkR4c/osVawznbrqSodz1
wBZEAO4DqVQ+cu/dqfDtFqhosKPLSuOkQrYvkerbA3LePzPoXaRa2nZdM42lcUi9G85iXYDGCmqG
UMzY8vY1Ni4YBvdOV0TJZz+MGr8+0UEaDKEFbpuljMEovhW2KcB8ybmtJJQ2Nmu/IOaAXnejodBX
ga2TkUjB2kowPtBUK3T+tBOaatkD/EHb7I0VvdMM8f75ZMf5sf2iAEcRuvOy82/+Sa1gzs2C2EFb
sfrIoe2iu8GiHiwXFCcZXcDB9ty5vnMSrPsuqxDOtBPQ6utZlnEDBMqNilmhwjnGXiqjckOtW1tS
Jxb5wPQwu9vp0G8s2ZaXCztIJr4SqLzeC2OYz0mZ4IkKYvHBmjwWXiDXXKBYrJwdgYmTyFqaFy/G
scItV32WXAIN/JLPJ51+UWXdWYUpDiNF4tSeoz+NnrDjHHIdGmobATGXgTlRAzZBNvFmhPIrGrn3
uN7pv/LeA3+JraL1jiokODwwLbnLVCBdRNSGiWnGbbRG761bGmo88eXMNnNR/fUS1japxKa8ORVo
nq/hTWbT4/s/ZQ6l+mL68IIQP5vGizisUDn98duqoeBSwZDRMEKZXZ7VDk1XiTbQP0a4RS6NY6Kt
iZTC04jSQKIqRs3koAUlQxXc1uMFwbOe4qeV0D0jYF1QOWwIVzNoXuvVr86BOFmi67Jg/0HXbsFf
b5Qc+9Gfeyc5yxake3TJnA1hndlgB5vu233X0Sbf6+Hf8RQe9Ve2eE4UtEmdJm2l+C8crYT5s//l
kccXQTxBMS7rJ5oMW51B97j/H6uTezOrvhNbA4ULRUElna83hPnohINntDxfZNlr3wel8Qk2t7AM
Z2bioIq1WVK5li5rZh/Bblk/HqVDErwUigq3siLEN0VK4LOeX0RnGxiDDkwXqZfddlmPJgdmJdbr
tkH69caK3OMEHoL8h9GR2OGw7luK2Wf2tBF87tuYifCUVtWZ26yjcLPWj/raxKRLrvQSWloYkpTN
fiF3Wcpm3BJuKuS759O631zZAI6GoQ3bLqIhUQYS9gszcy5+oJ5P/mBbu8Pv4qtESkPzI6KBiN+m
4ol9VSxGSTrbc3wNLXFu0DD8dQYeuCf0+qPUUKfO5gQ4AkL4DrFDV2bqM+wojKMsjLM7sv0crvdN
jwTsRbPCB1+1qYIwwmBKMODPzyEXcOifiI1le49vp2h/7R04bASxqNPDmrMgrtcdgGddTuLEPhJr
A44R6XL9x9liNUWie75SOB57G6v5lUeoCs6A8Iynru8Cxb9dxNkOEiNSW9kJIOu+2TqmkRRhxkGB
gEahYExCOVljEdoy27ouPhnnOSFSxHEZAn/SvWudaOMxjls96zoPolZ5oaNC3OO0LydAOd3AhPQ6
jIX5325xPbZdKRbDYK0Ds0U0WKmaGOatrqY+vuSE/nAc+5IEfFpSW1Vfo6CGziT6MHk5Kpm6D9d/
seNvUcBw1/0DEA0L+0+/49wx2pRJk6HPkZVDgGznPDR77EYp1mfKCZUPKPX/AvmE2H6YY2PYdw0w
vd0Rq/xoyojgAdWbBbjTwhO2ngosimPhsuPizgP4f5fIoUCIcFKW0uS2VySN9b22hbwhoz3pkPr/
ArAc4ZSGfWXHbf2X7TZR/pXyg3h1FgEBvBUwrPQ772uQI+D0OyILjf00hyT/6NY1WEkQDNxo436+
8LchJtc7VmK69TFfiGuLaAILn/Y03YR3kqblbnFm/qS/XZ1mMVF1XKAGSKvqp4l0AFyyDSQ2wGhF
ZEwAoV/q0hQyR3H4IgxZ9MTKJcSHUXnz6I+193F8VFGz5dn/qE6nBoVd8ROCqucHV8hakkbPKnw8
FL25QS6WPpeJcQEmuDp03ZXMZLHDzhjxmkNxqDdQPpOg5OelHvYt8w5d1JSqG1kxO2+KFGPhlQcL
+6pKWxjIQ1roYXjqg/Ci/oawU7ArieLYoQaUH0j8uxH+ORkpXVqyYLY4hC4Zdao+Wj3SFP+iohno
b9Y6X+m54dzbhMi7akkE58ho3+R90GQB/t8KpTXudIifZMBLlM32n/d4mejlz1YtLZibC0Cyrsn5
HU7BjQVPJfkGoondEPS/Ko+9TrubfeY/nE17uE/L6gdJ7k9LVF0BW/aqWzpV/r8iP8yOauU7H+0O
ErUPDJ+Dyo++lCwCKz9d6PRTwJcfveQla5V32vNMfQbgnrOdYiVzga7u/pvSduRseeICQZkElgy0
VqtyI6hkoifYtJHAIX400KBRmD7eqdbwTVBjuLn6KK01TgWo+P84EkbPGBvecT01CLPHoDnqoKsG
rgdXNnW0V3AMSBnJUSA3buWbG5QgY3kr8Jz9irGDpCeyf+Nrq+xnSoyggFm40E4kIzMpNlVa1YkA
AmN6BIwlO1DoQeJU1Ap7ZK29bz1jI9hzl6hQKWdunTouF1ettZOZtfsan8NqbgGwK/8e5T3alzke
6t5aJFbGemR1bjyDH0AvrxNCa2oXEw0VgxSlUeLNVbcPLIcfVXoqKbYSFKsWi8FVlWu9a0ilsRnh
v2xIDndapoj4WsNczUlq6eayJake6LtQflLMK/5letyNSxe2g+GE3oJxDetcNK5uFNL99UWvTwya
HaY+JastJspRqJ7ZwzrR8IzcOQ/HisRbOkiy2KOOZSvdCgt7yrfzHDe1p5zBRrlamFbAz63wlCnA
s11nYJC4mPImot/QICc+W86pCFGLYLDTiVrrI1VC+KX4j0lUN8t3Ab/EqXgBz9l3ywAfzS3NSFVf
H9T1mDdn9hIKYa6OzIiB+S+vb1CYcdyx6Qbi+gY6WirAcw1XuPZyGm3f8glOsisyWPs97w+DYzuh
ULHmNEHcHzATzdYozir2EctI6YAsoNDvGDrKqBSEpFFnfCyEHxTobVbyKmRlGryB5YJHktI85A1W
PSg6rhxz5ynsOSdWjpotqrr5CxdAkUAaV2taKZUJvALo3THLDJr90YwoexbW1B6yGF7W3w4ybFkY
tAL+eVa+j+xPsyim8WePSPKXxzYuVf+DEP6cQCDvUQUZo3F2WUDDGN3w20TtQE7S1jzScCOYjzoz
kZBnGI2wT2W560cq+gnwf8O4M1557JWcUIKw18zPV9itZjsGBZcNQIC6wrbBKy0fc2SlOROkh8ws
C6umZ4MOSERGKDJexWaVii6KpslE6EH1FM1e1Dv3vSD0PquiQeqAwxYDWxixcDXLudg49LX5vh0Q
U2jJQZi/fPTIZ0Nsxgntb1aIdlxJ00PLRVtmDYKYXt+Wco9dPmdAau0VClMGzEB/hFkdqLOr6X/O
gH6WIkzmdxIsGoy2m/VsJGqZBS9pOMVmyTarkVebuVOpOd2ndZgDmbZBETSUWuKzVE0QdN9reB/z
ZyhlSZTtWFDns9Yxnm5eGfyHqKjC5KxFv9+n1EKsGJEzwZu8N1p0Tqpq8JCPZwYfdqXQK+rhdCth
VQLatP3bMfEhuuFvSH+XHYJWJHfnxcC4b9hBpH7qlhEBJVMkKezRzDIfh6nLje4Q9fmb3+eOyhOp
5J0ZZJyuSRrpB4GhCKgKSy0oxk/ltstjc+MWqbi27cucE4KDgo3BDvBwjpVTv8CgEtrKRmSVJreb
odbEFDeVyM+wVJs/1FVuNC8k2n9Q7qgbkt95lzsvoIEFGbiv69LLQ/jEzuaddHcvyKvxIxsIT0jB
31cCporxuedZEMvA7BuLMhEJ0zIfU817oT8F0mNi2Z//597aVTl7zdj6iyGRxIPClIColzVHRDEh
W175B5eXAx/lt7W1aojyIEDA/flTwEQUAp6+VkVtAJFRuxm34A90gxY2IIMGn/nPRUyvbezh9RSJ
8RACssVQ9Xcs91xkCtGRIxnPPfaDZzfASZ4sEjjCHq6zjBDGG0Q38c2OozaU5Z5g3AvXAMGkNHkQ
46nYP6WV+vvGCZ7Z+JUcHwQzPhFPynvTFCwz7l5LIFMZO/sp1p7wcO1FTVdIRxpkDFKPTK4TsB+3
HmZHU1CHarslbSEofgC/AZ/DGQrURw8bYj2ZHuDDMbjlyANJAMSjQaY2OS+C5kIvXTF0+rk8/7V7
6HN/Mx8sogKZUV3VVstnGRMG3hKg1IMDWYWVzeN652ANA+25UwgKZssTIgW8e2qIpN3u2HN5ikBI
bu1Rhbs2XFH/B6fOCe8L/H84ftrVOc4oIs/X2GH6DKo5P75o0mEAM7vgQtC7RqvK5MScvGMU2jgV
7arZtgx2o9Crni1u5iBcnox+KczIauEUsl3qgozM/l16seaNLQkiEDgFHW7plMfeXRAc42ml5D9C
IXs89XOQ+5MGGJyDDOT7DxBSfFrx0721VyHajJxy4D8dC45y3+/oQfFhkojuh33R+Rxq0RjHHzNW
mqf+NQcR6z/QpakxaxhrINTtSUcPb7qBhrAs3OKoaG7oP4lGCac+UIjlR1kPUAvD/AW0DG6Wbnqc
5vtpCGl3z5YcRZAmfI3O/0lY9IXhMcon3O1sW+K2pNaNb7fvSKUS3uBHc6xKwOkyfqBnvYIHPnyE
21UoAIAfKmADIK+BPMiP3/3KZvN7CPH0WY99q2OTXd0pQ9ETXPWRu24/V9hah3icG2f0Fj+catCe
AsG/Zl2BTQuSI2JkL7mPPqUPLMt7BsX8Ac8pCHex+/tQ9eANjUGskeNw4lXPn+1B84X/1PkVWby8
R+NLTR3pUiTEHyc9JnssCzzlcskWJl0LDVzvSwQOrMocTAFMZkmaBTyL2C0ZMQhm5K3E0C6TATax
UiMF3YQ0mwParkN78Za1/4qgV9TuU8O0tfKVLNt/8eYxi3N5SR6Ku5J0yIwQ8DWQclRBwWPHzS9B
1J+gO/pGHBZ9xiUM5CfiiXlIWVkTgpA2+5wEGd/IXrIZ0+QY6ykByXWFiJZEJ7PaGlUzjIYeGSu4
gvqtwzMDhcOtJ12hoKlAS7wJYss5aSq8kExaQFlOVwJkIdxflEQ9O+bPZjBGeiSTzUbMGCxDgZcU
N+TMbPtw54hr5a3kYtseBC9d79fKerHI2UeFTQJHNqvRsXrcMFvbfGOzETb6MKfO4ziJYSStdb2T
3W6ScaIHXY57Z/RTazegQmHqqqdFDZSR4T1FCxECxepfTW4PMslFI5NL7LCoM5nPEc1WnniqvS9A
0npxeIzqaqQ2RBikl8YwlB/ag4FvDTV/vs0niAPFR9/zUvnGO3pdXRoQ2iaWnu7cqkMcMTVMPufW
qzPtWeOMqC4QyYNk3/1+rTjVsU8YZzBjsHzPu9diCv5yHTZswSB8ArDCrqD7/urNtho6mVIbJJWT
oJM7OEynF/wJ5MReLw7iQRpDeBtzGjPSNTxFNT8rAIw+b4OCSUVgFsIJ4BPUAOr+Vvfy7NY+gR5E
zJl5aHFtNFkh/s9sxTQjHk3SyQ6pgUbmG7efG9VkSaVsH2XIUMYMaFesHDUVrEqqkeZnM0MZD7W1
m8FhWR1RjDzcVIDo1r2QkuJwbU1KmOKDA0/NWgOxlawHjj/RI38NIexWB8NC8uvFpkPQVgY9zMha
bVhvTPxKE87vX/aCXhjRvCzQWIYagpFr4e/buwie0eaAwNr8qYF34O2kPV2RwPzbsOZ2xnN8xMUx
6jC9C10oybhMz+lMktx4gz/Z2iuC7ZRhB0z84yQ+MkXnjissamIV2FMR9EVcL57PDINBUxG0kdEJ
YIptW2BJ9az4EcqXxVC3aQkvIyTzD1GXo621ijI/W7BOYEcn2+Um7YfKKakb+LDTN/HPiwlUxiFQ
fm/ZfnljI/2bQRmj9eFVLlug1Y1McakDLUMQYyPNUZ07ycVfP8EEo8UfP3QumsCRbv8y9VPR2rXU
9mRBorIiIbN9do05oNmf4pYTxXHXNVj4LGkJHKsFp3ZpCZqP9rrSV7N4iLla36WwRpisGN95mae7
7swWAFpVDqxq6LTFLcP+mkNatrj7zfDjcGLZcyboigg3/SRRB2na9u5OB+yIRqbQM6jXKkCRjG39
B0oGCZjKuVywS3WPAOnFPSw3w/gq4PAbQa/AZG1nQ+5CltVzQqwXGZWSLgMX5IzdIcMp/QkuRr7O
r3fcTPyYhbTzj3UTM5UpnruRqtMmgyuT4RrgP1XX1LxAK5zVe2JOLoYauYV9uZqpUGtMNSioB9V5
MZfOymnyOemwxt5yDo5q9619xiBGih9aV3O34Q3prEnNf9XANQfb/UfmQ/0uyNkocGzONtx8/smg
pMc3rrVTKs0sFZ6P7SkKjssuiId5OyynV8wKVyomDjbos4j9iQt3SPViO1r4YbTR8DWd3EkhJgsc
cez8JmEEvs1l5JFYmsyclrpOvi8zGtrMF8xl4x3kRpfnwkcvHyODrhw3BSDEoYbbn6ywrbaAYYrS
l+yxpiAs8Gv/jGvgD4OBCs94pLKQyw7KB804yboTJFSQFVcMH5zQwXRdjFfggnk/YSdqpGPQrejr
dSgjsjp3VuY58WljeFUeAHQ4CPsjyR+DgxJjV7gO7Ts1FLffwfzpCMLKc9mg9J71WuLiMe3oiBoZ
xsaQiNUIKCMNzsSOOBehiy66p1AHnAZm1UP4GA4C2w5fnwhGYd9feFIEiMCMz7SkS42O1xhiDraH
CZiEtcfYCEn7/miWGAX9PCMRuRUYASeFyC9twYgxRAMXqvgq2S77fZfmjApp50EOlm/8/QMQ904D
mj8H18xzfOtXknYfQbEy1PZFORvykY7Sva13N0YvcNWPGU12yRgy3ADVts8xljqYFtVowoGsXdVU
EPgMab4u/A0Vjf7IkdlU8u1+hEoJZuesYi93q7nLArIktUqoIw8mz/gQ9k+Ld02fjx5FMcCEBFVV
n2Y5Us0MT45ANICoX3/lW03T4SftYO2wdUBPX8KcYehIdRKces/kJzS+P5IzY4joh1XhoZboeZ5+
uuDwIwgEkWdoNJbkYAINB6HSf+ntIe67dDYgRNUeQbnZC9xhyzbGbQi9PCObt9XdL1AE3b3f0W9W
vQiRKBly52svbbcoAMw7FCJfGhvxj63XILg29KQbLX5D3EbgP1hZlOWR1DlrpPRyH94x+ZFd93Y+
7s0O01rBPCNvJ0MtjYpvH1qXRALhqhwbvN2OrkHK0IHA/hFhSMEI4KRW7sZ1aTcwH/7VaFAX+YKc
jX6jraFnmzwgQenXzbAg3ezogTvt6A66hgzXmjCBNiPcStNZ8MKNfSuW2UwbEbkAU0nF/kN5Db09
ORYWMU/gqQcsMsg+Erk5QcLtMjQHuj2cUUnHvPe8QemUCFWYro53PN7gKgHN/tpUWbR34TQTqMqL
5RnYFfUKU/sLxgw3d6YzqftxqRrYnaHRX7708AAbZth2SrIF+63bE+s9R8P+hIxJ/ZKZjl9lwWml
kl3JB39LvxI7FVxkCExiMIWYMLadPYntz+pVHOonGVjvlBnVXSEjye6CFlT7brzDV4TxJQsWIS39
CFfprK0i4dAI5k5Zr+c7WGFUc2pHUJLasXxa4FvMADJW6a7oKI3kyQWdRvsrmPeKlSKpVUUP7eEu
uHYPloEm+tEeKdXx4hxB+WRKkysj5fCj8EyvFlABT3pOQAyvgKeU+ty/TdCaKJm5+UGZtDtk6+5J
AP1AyQibSd1u9bB2qcwXmtzEL6mWTspoLU3YOvbKEdA3I8yKKG5go4hCSquNJD+WR8jDbttAe66u
s9YRr6hcSkyOGixR+mN4raR1PeINMtnWShqZYnO7Iw8yn7DufDmvk9A/iIlcou3VNcbo7gggP3T+
bGoX+gsnadrCaRoPSlmucAE2gGVF3KlUTOPfjXbRTjcSLot1moqMJxphpN3O6LM+WsHb7w8UAAAY
z3f1jkubGNWpPh2XpmIMtVzWKl2E427Wx4tbWtXQaq5J65vmqcjKoEOJg7F3RvwyBVif9joRSqW/
hcUZiEyI0d3NC7NHn5BjfkkTzBUk6NXz4xguTtVxDXhSMf28f2mlry7MJIv5Ncm1KTwLw29cS8Ux
sA8yVjEuDcR8WPTecEJWZl/kzCPpN8vYCjfEcarYfHeVYXHvwFv96Qn4QMys2d74iOehJtjKKw86
yCuH6mj6/LHo01+Zd3GF9W0dgKGYufX9LIdzJVYDLcXv5vKuDwZQ1GqIqY3atfevh8uHCqxEchMK
yeCoTVGNDNIcd9N/9zgujUVhiaQxHELEEzrv3QOyI/BlkxqJ3zgz+/itOhVuDKA+BbW0nlKuJb5l
BBBUPeJf1DdU6WCt4AwbZU6TMoBY6P/ijecy4lzEuxycN92qgMUw1P8AMSMGNpZu6hsyoVUGEJuK
Zq+sdk1PRWO6p/8yWIS29XOp5ECT36CbQSoQ7eMS1ZGJtGl5VHmk6ofv44XPreBN9gLg6DV0N0pe
+4+Keel0lkv1/9cqc9yyE3iKtS7M2g640UQGT4JtoXcxYkZqfsIRavPsP73VmpbhYYGksa1Cf6Ou
Cz5nsWKCa/rU0W8ChATWOHk6vkrkHqoHMDrb27IuwXg2Qv2YmGTB85kCs38JQE52o7y3dAgUBpmw
Ur/wb8bwYaG7WAoxAjA05942yoWiSxTlWdMErrwhCSoUUieTACilS1yAySuncZKlitcPp7OLDWnQ
xwplkbfl5w+qcrPfgWSn9irsObW/hJBeP8aVfkp1qxCCWs0Sz6MkUJQdrai0WRfbQPHq2btqRpCq
iQUkq+06D2mA4osysKr1NK6ad0PjzcjiZyK7VoMkeOIQ0ecCcCG5YEh0j1UTzumsaWE2WkMpbAzz
/C/0caVqTSYiNHTtao77dzFIl8rF2xbIjyX3oPfT72haira64EKhUT+RXoaii9+eJI66VtbFpb9c
gwrZQysNhl7RxhTqppxBxPevvvbmyFj4e6QtM2oaZYRUK2GQH2lr3ICvwpDB8pMpkCcjN82pS69E
8bzwIS2FQb1GbN8SDUvg8skBlwIVKGBcwZvSpk8bPS1pcbH3UuY8UyGKEMeM26nqJc3ltKK58pzx
bjVOF5ny/5fNoaOgveEmxavQvcMjspXC4/MEJN27aW/e9KD1uNPQhlG94BRMZJOGrsJcjIu++/Px
gbA8dU/pq5L0iEd0BPRwjOk5UFsi2f/YAKtfNOCepjY8j2hyRaZ7jMMk+DRDnhm8uYjxDJpkGJ1V
REamk4yWdR7428kJ76/uuzGimHh3b0bnSmifo5H3yLO6AgcDONPrckMT1cRG3jiHkZoPOOssTbfz
rsv2QjgloNLmJifUCUfgbcatK6WYn6fXv5t1UPGZWyIyDGwMrGU9HwYaiPEozWPP/lNkpInuvRJc
Lk8bSeIttz0KtlZ8P7Z4gwCZRKpQu8Qg5njsDTaWzw+EFRpVXBLYIXAtPQ4ncohl6jnCW7TkZUrQ
1ymQ0qPYijDfkOFqnvg6+nF6kUzmvc8oMnQkaucO6sg1HEZSJ9K9ekcnHhbfo/emQ+uijt48dTg8
0jwyFMWHVCXOtZ5c8TD+PRmvg6as+KzW7KjJ1751zhw721+hR+t1OAuTuZyo5nbKhtCzXhQ+tLvq
ZuLuGFe1GbZGiCaI1xbXeFNUVKOykHJGnh9F97YvRo/R2Juqi1gQI+yS4vcAq3Pl0B1VxkD4tngO
Z+GqZzChfIdEPUUCNrIN8v9pR2m8eC+CIgk/xhgIVTIKUSFOInetbefozfDcfdVMbx4pwqvLOmy6
pLO0LSIm9VTxyCJRSYsXe6qhdX7avFne4WQ3a77rdE3/gaKcED9R3mnPaiPNpHzS1h2Q3/TEMypu
23cSQhbEJuoJLqpt53Zw7i18Lu191vDmnUBc0ngCPUO78sDwpajV9beXMk1kwdyMv1wWTy6Gageh
yDDIzjM7KF6UFXDCAykqJ85wqxtRfLRoSCIi/Rd5MNrkfAF+1+eJN1eExAh2OCFVF+ol5hcvaYgy
f7zsLEGhcOqXCksDIuSU3+cp3KIJiLuEkTpvLq9mw0kh0sAIuDpBA/JNW8cshjGpvBkpEf2o4sSk
QsQIoYKdupOCYvJ3ki9w8AZSOAp9QhkJXCsyrbGaSWoXoZ8JJEBadRd5fe2A8bt0/GaoTYeCyJGl
R0ZrLgo/vomDwX1ocUeTC6rAPTc0NfIjcFzIhgxfF0EAX1i3TRfTXx9CUAs+LlOGR/WDVyNNioWp
Gi6ju6Gt/R9WmRoKGuBPNA3zcnVT0mSwBtpg8h988FEJ03I216g7wcxRY2ZyiU20O+eSJgR8rOp7
I1BFHiI+a6WvzAqbIPvncD8DSwSeHExgR6ZADDCu77wZzKd0IhrkP/Kw4kT1KIxK8k6xWlvW5S+4
HA85HYMY28tVCAgeDXv0C4QkfhL/B8uvwGXum0cwBdqaYeXfmBNEHh3bMfPGYUxsXJ08rI3MPC/z
vdadbYBxCaQvFJE3RwKAc4EGLYeMjMgsB32VV2FW2lv2VLsO01ffZLIDB0Ri+QQayaXMuf3gFlMb
lH0id9tTnHF0hD26yVKegiYPJVwC6jBnQ64ORLYZ1+Kg3LMvZHPD8YPFD3BsS0UCN4k13tMCLt29
gvuIVKD74aG0WNkbfWoO2tGzje4RgCxBRgdpP2Q+CDBLVqo7Ri4+zi0j6PIYeMrOV6MnxirD3Vdq
BbENz4Xbti2Rj/YXSBrb8CiRZKEhY0cp7AxbF2mlPqRKaM6VRFp+CL5cyEfX9AHmiyKad4w4HbLa
2c51mTLQkIrjyA3iWPSOYxg9WW6ogeyg9s8vvbB0Wo9eSMhbKjrJKoGGWO88Z4QAXjtnksgt64l7
QBaRv8Oj7nQVTqm65zbvsd+VN/iPLfh1Kn709aP+dOj5Jtrc1sAQONGfvkIEvNClM64AGAMRFDwA
0RAOARQZrxfTn8AlRuIkVpIkKgQBQ2ajug2W9IX0HSMgexcFMrk/hr4SejmO8IsqmT/OUVbgaoP0
bAnoXMgBJ+JdgrlOj8w4SjNMisg586TwRWCUY4NiSfyCCAz0Nc94weahPve1l7pSWMUzaAgibic1
oSNGgyLUYKp7PLMpJ4TJ9kHB/qgGf3lWiSUKo2UD7iGp7MtKhixnN5rxLayERqwQSir4Z4ZivRy/
eSIJODOxbIuw3zshU/Re/0l+1CGIZwp/CWAJDYQebl3luDMd34ALf7gg/wShT0rZLjq4Bwy6TgZu
Ihqs6CIz1Xx4d8kmtpSaNcc0wSHakOkrrldt+wwYAWXiI+ymmCMGaNXKtGUboeaK/pe6ly9oQk+1
GOL33jsp/fjgSU4HQtXrjGtHDU8/+IsdLkxC4Ycw8i+4JF7CCDuqQfFQxaQBM8LYysMfyyNhrmDi
fMqSLz5tQqHczIz+pak8QL0LKe+C2yd0JN21XZ/wjjwyX2De2xsGa2T1tSp64KoBV4DUoZnBV3Md
w3NlytciD1pmjDHK9XcArhAwjhC7VI37QR+qR1bGQRO1wf4mbvKmR/l+J2zEXScVNZzl36SFUqtH
X2LtfbnX51IRui1CzfpFKJi9R4QHis/0N7u2qNtaNUFh2MRVu884tms/Tl7VOrRU5M/qZrhKIen9
PQL46HnvzhqocICGSk7ZCifj6S2gckAeyhVgDwu76rM6ISyqeNrOv0Qd3/nqKECv6g51Xj2CWeXu
oLj8o7X9mzCMiLCpCqJHaU60j2NVNCJrzzooTOOTUvp1mw2L5/URTCjDW8ZYnf8ZHy5wSBEm6aci
1OKqemCbrQMZrIyH4mwOLQtVNlbdbrx2IyexXR76PF4lTXZlFzXH3MFnILf7iTlTOiAp+sNOdDUm
zsVfXOO+qpXL3Hy3sgjYcJizr4KOkhJOCkLTYcz3qnTF6ymbi1yuptspy9yp018yO4GqFsrxTH4y
jlZGy5FDfqJGImAKXMWTGTLXgqzUcGq2cBJI/2SqqS847LtZcjVsTRCVPSI+HLIw6v3GSwQYUND0
IMVjr/CQV6M22b3l+EmI/qC9ezOWySiB734xbzBNi0FvvQZp06cS6FZSfrjBOi1H4N/4uk73zzzy
tpaH6hNKStUJOkJRhmbFoN1fJ8VUOSgsqVBICk366VpycMq+cZ56AcYZqE0/MN0dV7TAkYrPDLm5
P4C6qRtJIm+Un1K4KK17pTtm5p+miBPKgLJ73yHMXLu9S6meYVD686afxE9xCjgE4hU6LJQ2nZBx
qtPzrJ0oudmgFasho26qkZzsdh5VJOzjdBde9+lkARdiod9LmfT/dBUSR3W4io/u8023JvZ//naS
T5ytK7ReEmOmScoQJYVtiAIHDko6S/mzpfeiX3g0XXZkhAV3QhZB9bYoaZmA/uCfPvZWT7pBce3C
hkt4TWtRcvwqDdmqk+yAz02PYwurvEzTMBFh+us/SC7MMrPPP8G1vbcl/TREIuNJ+gzQ1erVbj8x
R0UL0g0edvfwbH9E2i1jLIOsVervq3SUHYybOdGbtt3G17XrVxMKwH228qLfUaLRvdEM9lbwKuQ4
IOliYtmgK/lmoNrOJ7DO4XyhK0oSmlU2XiFdt8XK/Juxk0ZmNZByRRqZm4ZPwoHKelXVojfej/TU
eNByYdbuoNLgzTizjiRip7RuAwN7KesiEk5dy05Q8DXrHOo9VCvWHo41pxEyG0fyrfFLrMq87Pc8
h/JjfKfjFGuTjxuCYFYUR9rEzwK4nzuhvde1Q1/ARdGgk36ZafLBYVmpOpOmNclfZ1q2Oaobbj5a
xplnDxXR7WoySkaxtIhEd5De6Pf32HmRXMLqbKQeVWkLtaIsCHptlXbD9JekigWxWlv4qYNdc+jN
RFECm0FA4eHxKGKfKgA1ggY6d/eT6oKHzwd5VQivKLTSmed9Mewnc+wM1pJ9TTSdnLwHYIyiYg29
VwEujPjkyBhfzERvbwLbXbBTMOcMvwqgL7cWLndR5nR+kXRmpIM3NzkgxHh/3RQjAN7buQ+dv+TZ
u+mKCmD5IJKkTh2tjHKQHAu9DaETOyrVe9l6VsQ/zJl85WXOyKoLLAk0Ar8I0muEm2CvZU5wgZHF
u5OQIKD7q16A+KsS8RK7nxOhpQOjd1B1dccmCBfbtrqrZ0OTFt0VgS9cKeH/7LYzGihAbDFnSRLm
eOgdULNp1La0nMLGy5oKbU3cCutLlsRSs/ylbDZPnGTlxSIsQF8cqzzTXj6SPoyFBD+R/UclR35l
HFmdu2xHxuKIRhZ7m/hJ1x3J3a5E/NS+lm71LPFE9tMcKJEjLHSyg/G6mU8MirvN0GGeBkqgxeTL
HVO0kCkafNdc9OqljYwkAf+G9mXGJ/7rUq+BzeSimefCVJthuzyH4GKGeq5qRRuny39duNND6w76
/onQu7Nxk6Gh2VjB3Q1lokaczQPpEHNc3EyjeIhBt09hxe5D/DZMRHU0uGCrfU01xDzLsvE+NbFK
2uVrAggDNEGh01l3rMB9jfxyReCeNiaHoJVtNzG7seuY1+xqmYKUth8LheeNfu6D+9x8k0fYSBG+
i2NAXyRoDsOLsm9fUjZn4YFnBkSf/YhWsbd0bn2Eo8bWHajP1/Ap133ZRzXkEFiEYQEr995JvomD
vo+zvyVr/o+O7hRa29/iHVVCFI+519rs5Af30PhR5swhULSjsy0OgRZvu5Q4Bv0clN9R5WqHFNc7
a1ek4cAIWtgoW0nakP7/kO7VWQ7HCZsGWCnZn9StFClnCQci9PCxxW6+rN5BxbLh8wcuc6kGdsqz
t/PZNg27onC0zwSmokP6rEqT902qLiMmjoxDlkB5WzZQ/ZS519RgHWAA83cZTpX/ZHuv5tnrXDWi
nIpqDvHFmMnyR0qzE+CrfbnUXyYjjkZqVz1cotIVZle/HJZD8Wdx4CA+G60q6mFh7POli00vdTbX
2kBjfn2HmjmeDFKG1Cy28d5afqvwEHzzPDWgpW0tgiJz+ShjWi//XNNqARTBIvq9mnAdgh0XK4CT
iKCcw4iQXmuzEy8wjxcF3ooUE8jy3lfzOM2y/8I6q1AOvTVrCglIXh4kx5nKIiY7kAGtCZxxuIOV
1+1sfp7IjRbhWisHXqCHzjER1uPx6rvB5LORX7L4K11wn0Z9EBjatnrCaoaPVky1wqSe2e4GlurF
Njdkyuylegt7Zbp0IpLklrN+9SqGJlay8Ko/QlDT75+YRwFUxI9zZO3qgd5YAWWpq3eLBxFQRcDp
wJbLmAjmPGTBtRDFuFrxshPX+S9GeCzoWX+5okh2oLQJk8U+OnT9d4GV2ufq/jJxiqjO2D9vMHXm
3KMwIkQaa17kVWNw/hhDnglwe0wWyFU0TZyTjO9O3YJ7DQtytaSSyv0E5yhsiuxePUiAS4RbFTi5
MMH2LvKuP4KUp63bxbb80EeWvTUvq4Q6ZBXU0lwjkNbOwTaVr5r6UDU7oAjhkJbpFBLRnj1RKWsa
q464ue8r8KnMxuaquDfVuxhHjxy3keYFWnJ+/YJ8sVuqo5Uf8/ldleHOxiUQGZsB/r0oriEalKgo
NAeWWJLXZQrEBFiufXBk5Ju1cKaIW+8F7NYpt+S/62VueS+PmTNQSK/fZ+lucx8lNg0M3hsEB8sC
D1u50vahpq1yRWyjoeHNr6cxl2niuE+GV2PjxYb4g1haEpyf4p98DdNAS5XfJ9uj8C+7b3civaY3
Euv3097yRHGoDGAlW2TAYdORdqHVtKD+OnxZ0pYybt89ltnbb1k/uUBH9upDo45O18BRM7wcuRwj
1OV7WW8Z3lCoMF8EMJHhwt7CxF79pA5546Remg6UUsrc/dj8YcCjT5raUiRZ7s1wmjHrCw2rBKdt
4wcGeTiR2/+EbHHF+Jo6Yp2ZKFUjYppfW5oh7sw5aqjUE4ocWTrqAC836e+E4nrV2K6G66WlO2Tt
QS03ILkjVVE8d6TK6qreP2JQtqVg/k0G30CVeTDw4vVK1gi6IFVO1EXG/7XUUom62ozAHLqbZudt
ars0Spy05zeqKawr6jSb82Y4AmorqCv6IMeELSKEJH5w3f3KbKeMceggFS9fPgEBeNWypYKEz0JK
oVJvkTUSDf2EfY/NbFTrtMzENo290PoPkWSlv79WENi1LxyD2cV7i/S+MllLlG4OHuoFwvpfyPLo
ivNyMqQO+KTO/E8FyRSk7AOMV7gif1AcuCJD2agSSLX1e2lO9ZR/nfX5iFwJLQlJBIrYplvaKpNc
66uEpRCL3h5UsWinEgfxA+gywt4TvJBQq4MI2RMdwwteDRQRFsyeBQqBDg8lnyrEqxNAyoy0q9Xq
gCLHLt107+84U4tEPO1yPQB3oJDgPVB6KeCi9aq3ZGrwNWXqjAj6NXepssaHN5vxPwTxRYzElyhQ
AJ3TgPB68D/4CoyjqLKGnxlZaVh3QonvZtWFH9UsDpJIGxhw7OUeEDAJLv0gYHdZU7FZsU4Dj+qP
9nW7kXl6yOXqu+MnpH77QE5nTxBb7e9gBm/7hzGKJbN95eO9D8WrT3+nANqZSc8Q54EFEq5kdCGv
4dui08Jn6gHyREhWHQ4Ul471lRpkfJHMDFWdpWpTn8PiAc3iCCnPtLPfgY9gMFCTBDtFvJMXfBJ+
K7n7yS10jPVvQz1CsS+VuvC9rSwO8rjaTYdyoEPacVs9TGLUmcPdsHEmkHqI+Kpb8odV0zgSaKyI
GcrwmPUE8/IljMul/Omqfv7/E0N8DPibLcpGX8UJwiStpT4OqFZ4CvBEZzn7C5R7uN1Ql/RSS6c+
hH8Ow17goVj8MX6J4fx1zdXWZG3OMFUZgYAgamBSKnf8gdGxcEJQ/qJS3M849elhxy36tlLU5rs3
TyxrECBTpnm/zVp79G/zRb23G2yN5tmVAJem6Mo+2i63MGVyQH4O0ssRjIwC+oeINNGnKa4OdWuT
8vS7Kt4JPH93Da3xHHjtZ4f/sRXiwahi/t8CKrv8Gs0Zd0PxWdkkcMKhV6Ykd6Ka9G8Y9mgAk3TP
TfdDxfdJKgC4ytRPwZbFtGS/TewMf/Ir7iT7N8UYaINB4xtwagJvjMD2Ocd6Rpl8V36Xym8c0sMn
3f7fvzNS5epTV4oJMWKLYzuDdAPrN8HWdfwXmy2/p/JhlfXw7IyPmoPCYSp+4SsLHakqKMZstjpL
TxudeCEk4owdfXByXfbi4l/3Xg5yFRdGwJdYFPVIw6vTvvbZq00K4oudlVWAjr4fYffbJYkYbXlw
yichFX/r+z/maGUyyNtspzAqJPtH+iWxmyxIQi5a3C6cYLmtWDXbCdjY+7okB3TE9vYHfise1CKE
TQWApd6pn6nRuyWxsqemYUaeHcz7gDbcvG/XjM+muMm/5zCU2qtFz5LxqZXmVOUF4MocZJpJPQZi
bADiUSI10Nx6kt/dBZsNLFqoavoGx9SQ/WYty+1TWpqv1syVUN0aGfGZ607KQvS3IZ6RjCvu948y
NknRUBE7qNYGD37SrxCdNIpvePmPRzpfNYNGJpG7EAexS96jnAORHa+pMpjsAzkskoWqWdvZEx+V
URaAZ6+7be8+RNd9uuIAr6AUhVWIYvc/tm0j2DB8MFQTtYNZPJvDfwy6RD+3fh3ZdJWf2qdNxyXv
cwTy5CatypjVXxv5RXJFsb1AKiNwp3sEMWSyMYjjwaZeHgXc/37lW5PWzZv7cVUU6cnCIu565v8t
XxbIhjng3WP4txpyuLHQhYE+8D7ilYk25qT8Q/8CQlmmoIgIqD1aJP1Q4Yf0Uzvwg466/OdxEVaK
bH8U8pSbgihSn18349B4xyhoxqvk+ETUs4+EztDqQsjL3r4AhbvmLggP5Y+CduTX/D+OlCFqBUlo
VXGDsvbG10vZohJ6cHdkwPw1gX8bmZFvOKZf3iPI7RETFdGbnrSlWG2WFXe63kc+Xxz/LdJtcVV4
EsbULLZkGxXP1OQpsAqcmzW2KgECAnZXYZCrWIJgz9sWFblH/OylGeMV4sj0r4eHlYU2aee3+Pm3
yIGTiDui1r/WIf/f6AgkzcpuCWAtAsXWHqzgoDgB3ovTxUNmJRgvZtq276dK4lLA7Xf6g4zVH9zg
QHC3wxeY3mBFKCpeXIQr/LO90GYH13hPF8cwQWex81VjbItj76+bR4KCXxi3ldglkk7rJaX8erch
AO8SHQfABGE9p2ReDAERL93mnrYDzccIpZ+Fd01GVDzBMrmU1QXzlv9GGzBw6tD3gIrXJ7UtEqHg
XQ6A4abC1e9TAl8/Erw41RmlcrJPOPMgvRqFqSmMrn32BijEs8gZDKXMvHDL6/1e/rbLTize9vBP
GqeB74rl2FBc+qKZyj+K/IKWDKrNyQHPCrOv6vKn6ckIp6Op5xS3rFAMt8C3rKjScLNRLhqbVtfj
y11v15OFigO0BlVikOuh0wx15BlbTIjVC9jAD7N13o8Z6nO/m+//mQq9dED7eIVBdYq3yr6oH4Cb
65rf4ddVolFGv6NbBJTsuqUgIl4VfXKp+vC3e3Bxwdt47yf9smtj7YgM+E7VWd3kecXk3NT46Ons
/c86ZKbL2agEUNbn2zi8u4nIMrdnpmTbNpHBjlpXWRJcBMS2ZewGi8C5/fNio/KemeiIxqjUSYEL
7aDwk3/h/dGUw73GB0lzAidmpUbFuXlD1+KRCXsgkQ0WH0yHOwgGv6lVWAFx0pdQHpVv4YAKg+LK
jnCIvpgSBjuZDb9QOFTaptw5vUFVDpVKCB3abZ8dMH57TOBH8juR1fidcNAofp3y9HAFktaUySDH
YZqd8OSZhKtj7/mFxOEQ/nyKZ8l5Jm+Pysqbr68U89S/yxJohKCWW3WvzyqfgiKkX3Wch9M+hqtk
zhAKs+03S4L8Hoc6hDEcfr8FYTj6HEnd5TXvuF7eFBWA/45ey8TckcuH9Zcs+Sl3PiL3fIzwCTvF
qMKH8mMeEYkXwNiCNg/yo+gia8Pg18ySfTJQr/FRhPDyUoxcjfdNh0U0RfRMYuWorMcq/DVwdQrJ
XxJf36FWMKLtZLs0fMYs3SfYybH8SkT5Q2lhjBlHAlwOzRoHSdoJtBCwg3yxBPId3ffwvLhjJ/rv
how6IJ4BIkwt/MpzuL85FhUkw9McJnFD/6mrbCzyi3Kdf32ouuaBg8uZEqnxg5/qRivM1nvlKg7G
XTebzyPp8EAJVIVXU++Qi3XYooe/s9HYdtMjVq/R2svUu9gLKeZMpkDfg863Qr7aJGodhZstN5WA
0DtdueB8zYuJozoo4G+qFcDYicZvDmHRCVPk36Ey+s/5tn1uTtcneMq+LoHqTNa0lJnWvPoBkztP
23E21vy0MZv1sHVk2f2UFQ/aF1ILb7gOYtB584sS7isXLMOkXMl7GBwwsnU88shcxAzPsLyRicNL
1qKVE8j0KMhpuTS7URERsz7ehDwJgi82O0HegBxxo2v6+Ex8RnYA1vkiC9l/orspm/xFw2ulIU4l
IrXoxiaVtt5u8bWCkQ1tfBEGAoPrdxOD/szuHaNw4zCLJ8FLt4R2wnerlkibl1qx3pvO/sxCjxPn
PwVWngQ+tog5sL21bISzmw5uVMO7Q1oKWJwfL3HJu8z+1SObuNGbZ6s1n+fTUgPNMYql8vbK6znX
9Mf42vC73jnE5nKoJ15jOkDV0lisqBee9s4jeJFNM86LGEo0CuL47cB4dZ/XNKkv6Rsigeagb5o1
1xhN0IuUGo5UxON+bxXDlR9t820yNWaqOYc+HQkycJhxvYkVMo4ZHWqdwXFuGXDo2yJo8mcz1muW
da/xYKuIYUbu8PS67a63PCKXaTOKbLwUipwJPKDw3Adv7PqDuwkSobNMZweuAim5SyeJAPDNmK9a
+cX9DVlPg9SBN/g5iCuzzdeCqFW+XC/Vc2vYCT0V3uc0t+7pwTaC8+385tpIB9NGZoyD1zMAUEYX
Ga1z66qrQe5TURR5S2IX1ipW+J+slr/GXYVSTLjGCB7c4IzaVJzadMPrawj8KtPu5sNHQRu0NzKq
5teNurApy9HkM6AYEbRz1/I5a13SQVlSbI+Fw52LgDcgH3rI/rv5q3ucSLP+tth3FcIIJCKHnXGX
RkIgVhD49iuFsOvbaYWAzAaeRadcYHNt5HCkayb7hUvU/cOeABiI8N3eMbiTycvuebeyCZD+9DxE
98RCOvJ54Km7wvN3yRibGp4nX6o0L0T9HpgKsRoDinNka6r5oAcVfiSzPphMz8kwwEMWvIwaWA4d
ce1CR0BlzagzSOogX127Tc2KHL/MTVZuFCoBfg3yyZXmpFHxMKnJGk6LOgWrvtaRwCC/Bd0F/VwP
Sp/5+qn9EiDJvDa0D1h9EJz6LsfmP4vJwVCFHF+B5mESuJnlNigc96H7que5ni4wydgiJ8yyf1Ma
Pl56+dq1CqVEk9RB8nQQqEcsgxSX/a7gQW0zpvEoYXIbJMpexYnNw7DYPdRQmhP05i8nSDPzlE9P
1smyCiqORPaR9H4tIKJAMEyqMi5yR+gJCuXOisNVEj+Vr6bf32Ugdr7zYT05QoiKocXvRGMnFcEa
maRpkdqkvy1tlDus5u6GhDbyb5LcI9hDyPPp37CUbGa5imlGQhj+MqiLJAiH50kNKt/64xHTt5nn
+120FAkSBHa9U0dwJ0T6oNaYf0CusBaPEXIoQ5XLtk3ydiVn2XXyxKoW0qNXvXZl2bdVhO1Rj9Gi
ZbB0B8kv23VCfJwhkzMZtdw1ZLMGXr7YTWwYAvgy6arOTbqh6b5t+sf01PxT8tQa5tiD577k/rrI
6lliK11pqIknhxWwnYClMXQbkMSzCl7ag34D7KylmeprlNC/SyJ+nAEi9y3WTfEKN7apTsaqOUCb
ZHrZfj6ed2S9rkDd7WgZESgAteqr/Ht0Ygc4rQygm7itRr5gpLq0wLChqBNkrAe6E38vi84vr+Li
Qq7qYvwJUS1kZlxe9G8xrz3lamrdj6ay2bWulFoW/UlgzKTbQQWWAzlUQ3IC22JrrnPPoM7P7q2e
qx34fFFgCl965LWNkfMubceJnmiCUdK8SclQdukamtW4IxhadvRazxw/eaHTi4akTyY2eimHzLw+
Ha0rYt0wj05iMirWVvLbCmJHDMJhV3NHcp1pTBHVeRi8GrUuRRnmAmemZZLTZqPXG7PycFImwlCP
WhFY3jsaRRdQYBIha1BZ5PCb6Ee/1ZkTkgjxASHo3ml58y6dAtwhqzS/NZMKcQmOgws193MQWJ05
fySp0PK/y80hvs89Ge8yalXWBK/uSKd+fP8FIsDyihtQJfVQR7zH2ul6lWn/8UzmeTE9I9se3ka5
foeu0x1lDCdknB9uqQEVuQ+Z6JvAda5v5KzP0IW8r3RlPaefFDnGMbh0XuiFekWXD3wIx+Jx/KyK
jjTUktr2Qhr6fNlmN8RmDJ7CYHXdTi7Oi/0iedlfMPwHXzbqG4lHez9tNBC6Or1KqK4V7ehO94h7
PBqa4c7vgUtyofQbSxiUHN8Yg5/1FKCb92JpEZ0QD7geC/5njl3tVSDT/UK35U0DaJkCVXR4rqLz
MLT+o0IenYI3+IWi3stGI+gIe0aw/0/97YIeIISbaGOBd/tRK33cD3eEW7LwWAoocmeqFjxaRLq6
LxMSFbhyhDrRZNcv9FN71mAgKytRpAGhtqhDtqh8TS0cyBDHhfPR1AnQPLJKQs3qnYo4io7dLRQf
DOMBo7aJWzD1l4nnuu19FMyVE+Ci6IICbRsePoH9dYin1cmhyatHd6XD5m08jk6rHI9m17FPnWW8
RJjKFbbHFbvIfqVOZnkQYzHfg2blN2362RH4cYLpb0jpwrLQ02LwtGyDE98TULD9YxbT4fBDHQ/S
t5auXbsVv+OI3KhB90XEzgHs7JTxD+g6TwajbfM3pF5msd8VuqhTUb6ATufXV0M4Trzu/6embT0o
dXHd8T9c01OvapXpYqzH8K+pSa+y7wF1/iJ5cjlfvtv8mCMbavXngDPX5KkxT+hPr4e+J7//I/fk
fR61BWwYFELCld9RRB+gN8raXb/vqZWADZg5V587J1DX+p7r124usSvRKLGVgjCfmrTc0F7Qu5/7
FCL81tPeh0tUWADgeI2UN2F+AvUfyARzNnwaV5ewY86b6UNjt+jKMsN8pCXzPRcYTcOCIyWQBX+b
nU8bQJZcIYOIUeXSLzJEgIBtF+dri7OPWcjZbaeB5oeUv5uV/CnTGE6l52/NOHLjhhvwPgHRkaai
aFNxhA/ixNSmOzQyXG1UAeBamO7v9/RH8d18U/OMscjGSG/HfI5AqIpWZcZQKc3R1DZ4ON4SiOkd
GkUq7xu8hAB4NNCLUE2+Wm3Z8yOlIfFxsBAjaC3Hxs592WBVcJZIbJa1tPysFULvKemOIoJ3HnaX
B7EvftWUVrVBOVMP5lfaT6s8l6UOELamOkQblJcvS8W2U4YuAx+D8lSZ/chENte4vWhppFI+3cnX
UZyU1Z48mPHvA/qUPqx6zdbRlxhc9WLd2l/WXMMmfr3LbTBykX2/L+Z0+nFR3mW00bIV5n7pdP3m
uaMQvt6lygRnf8LayU7QCZweTpCYSG2+ZZy5i9JvPdPBKNRZOhUcOQ/etqbCp9Dx3iMsS8oNjljs
hqRf+UYJwwRagv/T5lX/1Px3GS9fn5tB1gysa9doHybRiSBH6RHXlzDrj+EG9HFU75EPfx0n5Y7l
V8mx/9+RyqkPOWhtiXcqSC14CpsrRwd1zI8cG6d7tnX5J9L6r3kkj7b8+rLSuxc2f1/uMk++2N71
RgFnUdM4v9+m4TiY2Dx5ePDZaax7ZZzF4eSoq6vzGK/0rEsbOLl7J2n85NeLJ/JYoKSSJ0hdCeqJ
Ugwv9caaMbUMlvrQ0JONWUgFmT/yOEx2rxcI/q9aqVDxtqRZ6h9aKLQ4+d6qIBu3FC8/rGI58bNn
sPh/ya2jd5qc52faLVGorzdSArOEIk1RmnjtJ9qWy8PMbfcEubbvyWIQbwKNZd1/fAzIFnH9QMiG
wcMnzbzfAfbtELkkaOUsUjouYbmcvrWnxRckIpaK3A6MAzHbU2WMj9UkJmFUzjxRMZ0iPjQ3TUHO
AOQUrjagMXnm6f3joUCGdxq3D5olHJ/8H8V+cveI29f6aLufMKYmvoEjpDbn4TiTgPcrjt3xwJnY
TSlHkdlccQvxRk+EnP0PMz63ALLSDppO+H1hX5snLCUxzxBDF5CNUdtD4MwCZfUpfJ0hmEMz+3DK
FQd/f5SEZ8wi5xnrComsorVNFWfsx+SiAUpCvK/ifIwOxkJ5FmsWl/Wm9IIWJXWS0vunSnM6gy5X
6WCy4E/o33ZFpC3B+hfG7lyuZ4w7BE4w/iAPyHAd8C9VF3ToLFaDEHuDh/JB/BYa3aB5vZprntqs
DulDD+bLPl7XLF9nDpE+Y9xLN8ZsAzzQqD9BTpp8V8+y1j1l4n1+/VtPPg1ghPRZtwdmFTqnuTQa
GdROoSt+7EEB3U5VS9ATveFAHbEgYCMECmkXrWK4VOT7TH3zpzt1npKZi5jejAL9eL6lK/ZyNCJG
iMK1+ZZ/nULa2FNi1BO7pqbOs64/w2xqJ8t2YzQmZudyD7Ff9rRV/naE2fm6/2srUDQ6F+RnGCxo
xYtxwYRZCO22TeWQJd3xKyHoZiDz5CgSHh4hY1FrJy9mC/uu6RTTZNOh9Zzp1YhqRyU7+lO6Dgmx
+RdmFp6crJYHb14sYZElP5L31AulUMFodGFbpxqlwJLmgXfmAzdUM5qLROMqQ1JwH6Cjlhvel+IG
gLPWZ6Cb9dTUFAxkmPHZe02TeXEFUbwDwu1WV1fPp9UA7AO3k1YLBPWGi0AYU7i8vIJHCOpnUIDI
BEOEc4WQJZtFD1s7FbuxREzxBH66FN6eoYCJCaeb+RgZLQvNiYZVriSQTnGQoS0sydGAViuyZigM
TkzFF4f640ksmLwZg4E49Let8w/TKWN3v6erhLmUxo0IbXDoZEtZCqF1eIP6zSm9uxfs90UXSYUL
4WJkhFdIL5aIADgXhhENk4em41nZZi2iZpwf37bdxrdJWkhE5aEQYUjgW+FVbESFr37okD/56Qtq
gtXtTlUUw97I50fUfe3Pmadvy66Nl2Vv+WjxkVeMmXQ/KN9Oix19h0Ra00GVZ1HDO7Id0OcFqwaX
vRGruncTOnVOhqhORa+UZpp09F5YO7/mR71LcW+5/nwpWNtSUpCnwl4C5aCQW7gfe74zbGrnfU9a
gYCx8/ZndCs5vqfaIpaDD7cnFtwneYJ8bvqQBa3tt9VBsF573LUbHXkbBPmcO72BLAMkgQYm9oF9
eR1U0bW3fcKDkSn5GTqN4VHF3Y/Vh9l6SZf2kaERnRwrAHg9TTMG/7FMzFby89+iCKOO/w0CSMaQ
lWnSAD/+tpDsc8hxzPiRnrXafx1Uyj+qIoghuYs9PaySOnvocw4Ps9zw1yKqbakFFtQRH0fcSGzx
mfEDLRvy2xL5giywgY4wL/6mVA3GnQnyWHf2TG8tOhtb21OW3pDuSnJ4xWTHHLnhQhikSgV6Q/7S
FbT6ReDi+ulaukKQeONfQ+Diqld3KuEvPCnGvCg69/11BwPK9gCo9JV2ATqJO/oLuUeZmC3ZdPQ9
B/cKyrLWpdyJU+CVjxG+eR769roKH3WHgPxa4ngwKTGK28Sz8KxSdIAhp3sCBR5yBP+n5Z07g9Ee
cOxuIm07ZRLD9r1aC5eXqXzwmsUTchGoq0xlqx+DmNet4m5Ux+Pd5FBoXe25BT1AIBinwRETsthg
MeNiBlDKE7l6aF1LuHRJ0eVGVLeMCBxAkhQcIrgNkI8IoS/ZhLvfOhIBeyktI9TDagw8YiUf5jZx
X9etRBuup79fU4LvOOcp4EwZtM2qgZAYqtvtCjOqJiCItgWxlSDgDtEYjgSQ6/exix5LCAnbNmT4
kk86Dl0tAiLQtm+CxZ5mU/LLL2qOCiunNIxAoKYh1Op2efS6P/XSl4uy1axmMfaFZQQi7y4K3fSB
6H3Jpl/44tQr3J+ij4yRv+kw4XHVw2UKYbVdVrZOM5arqa0J9VV3dtQ8vjK1ADN6ECaVTO8zuU4W
sV9RbqxDgXLBy8A9jBt59uhnPEnIY2tLv52/yNKYOb/rrdBL/2Hgj7VPmRL4BLlKNUUgM3ETijU2
lLzrqKpop/FvymMq4TF//FyXzIn6eg+ans3ZuxtDg6ArHQhXP+Ban8HD1grrtzook2jxS0YJXYLV
5X9Ee/fZoFJfz/XTzXb0Hg1HaqP6+NAxATheSYsvnNYI9wc8b/Pi9DfXEYwi+tpA+NXoUnVsmgm7
IxAIQoQwmd5ZxS1fYL7D1X9RKOwRLpfgLtQws/fqdetza+Zclm3QAsZ64pvxAsdV+OohtPED6Q5k
RRuWJzwizOZroZvogPvTvLy/oTRwQAkfty8UIp2Zz8WN9Rxn26NP1KqVbvcgOCUphxEyQIwKoK3o
nrgdDvGsvhdD/P1pNpnqRvcaIreCXN3mluNSqq6piGZ+vq5ttBiT7X+Ba22WYNe05RP46znCeJVh
rjid9ewqNP5tInjPenz+GDLUbn6MYlGz1n4E/GOuy9HHIJ0+HSln6GcvxLK1DbYC7mM33r6DwE/B
rtKwOvRQUkEpERFSnjNZi09uv+ElXS/FdHlu5RIMY92IIYru4usnjNL0Q8o3rcL7j9OXsyF3g3h7
jBnNZOJld0nmUNhKnpa+xautVDhVtMtRrfwgu1oLtfI=
`pragma protect end_protected
