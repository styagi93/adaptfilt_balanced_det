// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
t42S8j6Y9MPyNFS5qMQHWs76iXGtZqIuXT1TarqM3yOaMLCNt3kh0H639WKGvayabb1PrQk9p+Tq
v0tH5BZdSfbThJycRh/X18CfcurJRLFubFrERkPqI8voePdcu6y/3ex8mpuMipkeHTICDuhGS6aZ
hTmRjEQXafdEUZqyo9P2glCesQptGURVVbOTvnNT6aEJSWYwjsgSXPoidO8hXsbIUAFL2TOTEn0A
9vbDM+W0VBVLVnnvpvrlbdJ49NJzjMdzyFlv6C5lJvtToSNTIcbjHveLEWhS0XKz9yRHlF73U0cv
N4JonvMcRutDXH71F7hEzXbTJUBCCi8Si7NjKg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24448)
8uOJDp4xhM1Msc1WFd8Q5Y0SJpVmjyVPzlhKUdD8JfjUCD578oGi8p1i7demJw3n2QiyTJIlw+OB
64XUIgudiVRjWFGe4hV1kdgNpWCJoeIsoxAtNEIASZL62CqmObLah0dMfAIXh0IZYYdQEdis4/5Y
59yI2mUx46Qhsz/MV4d+qn2EwCHig1mmB6PQCjZg3pbypYgsPWNPIEjFvX7ZPyxpRmVk8E8qN4Gb
U80YFgfkmiEUaoD/I7FDf93/0hzzaPbbO2YoTt4ITzAJoRXeVT7KNLobCBvzLQdsFIzGLjlyA8d+
0JH6Er5mtGdIigDVwIOiXgS3+cVC1OQjeVyZiAaEQOkVDfmK5OfdYHiTBLmV07LPjHW7lLvAXGz0
VOW9qAR9f1ZpiipMzDhmNA/Pruy5G5epI4EB93zrK1kcKLi5LAZPdbitMEefIWiqdR5OiInOVCSx
CtQZob3j+RHG9OVTgO+M1DcWc1K5kIbljigz2yHjhdZ0XG3yXnl2BOP4834i4GuiUD/cP0lNvBVX
fvm5izeNqdpCecaDj/WueU5BcmISnyToHNmEeBPJAT7S/Bff/mo/PkBkTjO87+fJbUkN/2bgkC2N
Mjs4UNwd6cc4OrU1/NgeW+uD2jL9bFbrIPbjshpsnwwUcDbs8dCwOa5eSZShDHX7av6/dpDt/wpU
RlP3UqU0jzlWaVh4LIUCQ737DMLp7Vrda2wmOAMVLgZ8l2R+2eT2FXhZ49w+sRmHOOO45adV+lrp
omSKeBztHVnGJzjvkYN/ely5ZIl5/uA0SdMUH2FcrJ1/R3aGokwhjDEQYp9MU7Grp9bh1Aul43GO
FkRG3oTf6nGKOhi04Vrp9vvU2TTqO2bq0+/54ClIzHeZ5UTGaXDTc/OECYtgL1vTrDG0lxoQdmsC
unqQUtrR/6CL590sTGFVRAsGcY4TiKkoHOaDSvQSu9b3VDt8PAjxWpDre07mFTJkGSxmObi4Sq92
UzIXYIdf1ygt2PKf9l4N9gHzxoybyPMG/jDXXmb6goAaes+A7uZ6Fs3c9BmeZKwXIXk/bQSDNNlp
j9s/J49qYtQD3YpyVD8qx7twTGPIaTwJzaskTUAvvXXoNvt0+N57m5+xA6dcP/U8aC17avQ/bluU
4vtNilyzR6n/tUFr9tUlGh00Wj9IrXdwBmLyvCEwOnwHE8djBYrIA7OHY57s3r4H1lwRipvlbi8N
p4b0WU7lKKEfkE/cKEH8SY44BEijO39/L0D1g7da/Zcj+a8e6deumc4QXL+E2xUm9NvNwOJ100Dr
oD4J+68D12FEmdoJzGs0a0PoCYJZCMIya5HOqdm+iw9V38OLr9192QM8kATSwZ+nCe/I0ffC3jji
Ak972qYkCEuKstGQjFU2h1p0CszcDTVjaajvxG+k3h3Ixym0kT96r9TtArYphIFNn+o+RRnoSvOo
9r9YZogHXch5SUCINAOuI9QeZETqR5OxidMssscLU6Vbu38pyiZpEXY6iNf2Dshn8XGjUJjDjUn6
B2dYmXplGLlX0PRCYvLM58zoDLW0X6ckva2JpxAlTlaqqBxzySAOjYT9iWLCFE3jIP8gcIAQSAkk
qxQvUzKtlyrirKYj1EUmf84mERiw+99raEEP+jOKfqPZvHqLrzKiLsQYbOl6aWYj07oVbMkbTJLV
ZWRwyRicCIJ6K0fHXIQJ2n5M+ZYrd3L/E07w/+mg+Nq2ckwCwMWOJel2QTwH7i1uy+sxOcaXH8/p
yMOXWd8UAwrwryHzsLT/Fe6q9liCGBgWrm7NTspk0hthlSX6Z6rdO4/zPVgDKkZ9KAXfelVkOZUM
XmgLP9AIyttBlL692BSUjldmbFvFvkkLWMPTFdjPkswuMff/BgbgKQEkKq/EU5mmK1dRT9cxKomT
h42brOGNap0dFexaUNIWJDpVHo9JGYajK51K17olXjl4utTBIFgz1h/9pubp39sGhB3pA4ZPrAd3
5IYr/ikFlPuoM2rOsPMIuBRKF/J/QJHS9kuEDr0jsCayD4igRyb30/UP9U/Mq8wHsitqU/KS+Ox8
FfzjiT+yQR+FyFApEohf+4OddajEugZF02vM7ZF6KyoZXltwSJkHMXoDTyDAzb4lVSo550WgpPOS
KKkbMfiFoADms0+GXL4/H5FqFOO7d8SMs4A5zXLaPd52q1e/zP8605HtMohHPwnu57gtAMEVwlb/
vL3+uysZDiYwnHc2H9/S9YR+RqNc7LCvUcnKdySi0hJUTnx96GzpSFJtG5ACWBQuvWKbt21qh1Cg
aeWPweceB9n73UdKjkV0AnD0IfCWt5rZNGTymF/YY/XlP118Aozns7DfboaWE3v3P4WRflcGubuU
yonjja8CPFLgxGNRbuKC87yzGh4iSSNq8SM7967s3LNVBTZ/IL9Cr5k1SmcFp5FD9gMzkhrzhWjY
HSogAt9Io4ItroQm6iHpb2dmM2dozcXAQYCyxARLtRK6qc0KrSpoXFkje3bBsjc2D+lOhTo6OfYC
TtC/ADzLBWYg0LPANqkbs/vwC4p+3CXLgAhIJXoglpWIQ5vHhZf7Y6+4BeE34PNgznjn2cqP9FVo
WczkjC2Phr3JmE0KLAkGeyKygNXl+libz+rHoSVy3d65A0FmO71ixrRZpM0YRiQK3nciTHgHM3JV
0s+JFWTucYmZIXrUpQE1K23aJlvib0KoD1dTdu9zaJuPEneFLu38sBLrz5gf6k1RYsXtc/U5uJve
zTZlsq0CgTL5bgfiKEOMs1Hu0/rnEpyzLbyC6vERFNoqVNEDGvwPogO+iJBHttvsTXQDZP6F5REw
whN+6x2IIzz9qz5eF3x1e7qjoV1vqloM58nGnGHgk2V+CGNxNirjdd07lc+4GPqFgIKp24YbfCDZ
Dknpe8wslijQORTUibn2PtfXSDUUBacXl/+zB2gqZdVfbJxTqP9QaIZ5WAtuK2/4APa2HrXGJgoZ
GQ0T/GEjjho9YSekizMuFMSHEE4rF9rBkz1JkjmqPfv7lF2N0atRkYJqEUAUidhfC+zzDrZk6mmY
R8IDlxX0QmDhtRoZqtQkDG9LgEOLXxd/PrEOctayecXlqH90ZTOPUYb9/j9dr2nHCpda/OCs+WFr
3K7PSJq1cb1C1yAdrd/zwq0hhnxh9bbFqUdjwwpnFVP6KLMOIoPXdlvSw0e0zeipzA4S8wM7bxTj
pf7exSP0Mxj7CjHkvxiEm8kTp2wCv3xkMYvwtJj0HtBu8EUxaWHqXcatcdLgEWi/1EIxMKby7V4s
Fws6GLrlCLQlsQPJrpJlBya95NpzNRGcgFGTSWj1D6fZBqdy6Ln8nTg0ozc9IB/6+pgj4vWpN25e
tQd5gzbIV88uCmVlaQ1I/+ReoRx9/mKEdZC196zpuXsRGAyBjBqhF6njsZqWmulk+HStE4AVgi+b
civhd2u3r1IIr8HX1YTVPFXqTowOr8eK4j8YQv1BqCUiabvF2iyuz4/sNpGq8O6wwOzn6lY66n9r
BjKYJk8qu+s9QfnahshZ1LyRX4qH27cZwsD+BLHinHzTrFqgsEbP8xj09m31N2SSjkqwpsGpIrL7
0Iq2HyX4vxbAXE0WX2wI74pKnhu0I6eS4CSRcAi69LgTlmGNiTqvAd/HmX2p5EaTwxS65kih2q9r
doKM4GbiZUKY9HWWhksyPkSo0QmV8bB4tILnLcUDPcXtxGHLrpJwj32IQ1KlG88ho5pVN1bwC/An
E4Md4ZrxNq5PfXYHmm9bHSJWFMlRzHYRz6uof3GfoyX/jALxrOd4X3snRvqrcwURH3FgRmjHNgqP
n4AabwsrF6Ev1gzg/HV44Ll9hv7RCeFeOOLYyLcww9ZEL23hqf819mYtPVMxIkM6PqWbXXhu6V6c
/ebjcuDBDfephOtUdW/5GVmHqW3GpE01qJCB4+9IfPZ6e2WSMLJSwPCeIoiuyVH8bAwTsk5ampVf
NBy4l7pY6wgvIle+OwffvAcLDGpqtlCrt8iPOrCamtOsNBxX1x2jYhwtz+B4m8PWPPwk1kCzkWui
KfTEuZDYGOF+C00qHKc+octspq0K6U45qvmOpfDhhARiVaUtNKPyHiHjHn6mzR0b1a5XNM79i7S1
vKLFPdWlGFVOJ+wSPuRLImaBUbK6VUep4Q/K9JW0RBguEVRLox2+OnCbJZPIYuA27CHng4HuYc2M
eSNYqkdtiNHs5EfQFkavN+A22vEmZ9h4v9PAsXIed82ZqPJ0FG6d9AdubSNPJqtglDv3eaha350Y
42nswZ6phEi7Q3UHGmmT4lGzGLVuy02gnJhn/gieGGN1F8Yoyq7w3HwwhbXDk5rf/B0+AgzobKBB
o90s0mmJznWb9L9sMqlb4GZqF6GvYW+uau/0Ft0OiR19W9ctMv3YaoodCU8lKtvWn8E4yrdE42d0
+t7rYQW8RCxb8oWV9D85WXEvfLi92Bbo2/apR3F18fi8JXzmMD2uDna+oxzr/gnzwiSmr7laZYhe
4NXoNhi8Y4QuEIgkLmtJvmPjm0pOg4bPSYD+cCvPMfac6ElPVe5lvwpd1UHU/Al8VfhPwCBXg6WK
fLinkPq9nTfrj42t9adBK+XtP7M94E1Ayk73aUzIunHV+3BjsVm8YSdJqoVaMTqJHbJbQ/EpJgZR
KTSRFLpZgOSXnM458s/+MFsQzvBj3n5ovSSgUxdPeWqW7koE9+5LQMHXFRYCq29IJvCv0QBanPiA
b3+sXc30IwuoxPPnsIEOELHra9UZ3yxvCoRaZLoDaN1uCZuwEOqzU8y/b98vn1WOgkM5nQYdrMf6
qvB851VuR/gJgBATUj4fesO4M7Y74LuCEgu3mT/Now2WdDdjdL+7rd3H2RfI+dLyiQLiqFQIgKB4
6m/Nc9xIxLWXf9uJIrosfwyn6U7sdqAN4LOUdLD1miZsijNcJgebr28CM77tozj/VIEdVpechHAJ
EHbjbI7AUjPa0cXITQPZpGN8t0FGHFKcTI9Y1p75Zmq5HSi26Nh5+dCQE5fb51YjNgbTQa02IVh5
YA6PJAjfG2ZUtM0oyC8U/p+b8Ytr2RE+d8+pKnR/3qsAKEE8ZqOqmW91khb7S9zea35QB+Mquxka
3qU1oR99ZZslCQXaGT3QU0N8knVKjtfO7t7T1+YEbTgFPLtjERRvsCQ/YP2ki+NhhypVKeycljwq
xYt6JDIsOMyca91hS3bN6Vrm1jypTtgBlthz0Q5VqIC53o6PnoC3Clsfs6di3d2siiFIQmQNRrf7
nsJ+jZ3teBA1ySl2WsYYWgU+Yl8DZjotOXcs/Ca2hmCy4hBysQRCuH50fCmtL7yXfvJmXAPfs2ou
JZtLVlxw32VviahEiTy6A90VOBNmkmPkExbNIJ/cYBbeUCIVwhnMCFcSjpPrIiJkznTYT43yPqCY
kITg2Os/KQjKQmQPbOx1SWelQcnrFjU1egFTpprUs58FkCbSBh5mDAD+/PDcBnJ/QKyTxXx312Eo
p4rfNQ9YxynMK4sks3Ejni3yPqD9ui+raDRI3MxgcdV1vGwk4K1uRye0ym15qYlhUo2BJYd3Q11k
njIOBEhh+z1nrg9PukL3EBY5/WCTgGZ6tdZCxTPSZMy1jajxaDdWRb4IUmcZOuZrfCQ5/GWwOChJ
soi/hqoPPdcbf09HwrdEq2T6EbU3AyZXN/ppZkZHAldCwYcMOgBGX/dnc90wh+KDmjrjyMFO7TiL
PT3YA2wElLC9FrHoDF3Kgzba37B+0W7yLE1E6NzrSL5pQ7bfO2qVWcnQFAcXicsIzdFm5GyQqDt9
P/VSViq1ODyj3uE8pBZTDDHu2dHkMoe+HdNDBZ0GzlVTBNQ8NzDp+4qnksWxx5IfpF7mKy34u4ZJ
R1OW0QDuYhEkMbPA6IiuTlRdq+FwzlIn8227kzUplnaFT8sDaBlN4dSeg34qI0CPh/Ca/ODTE8Xr
MZdHyZ5VXEHm71f4CdNI6WT5SEuaOpyHiu219/RO7nKpVhFt9WtXRJEtwJwvRCfBA4nhSYRTUqST
zbfuGLd7c4gK9l0QMxffdubsxlTznnq2YhIHAIa8lqCqh83NhAuut0c6DA3ZpHAKZx3U1Y+KVxR8
OQhqh2lXUoCfDPEZmqsq1F7pTqADyQA5iNxNjE8Ekk8o4KKErFMOEE9VAk6fbQYkKoPQusI5XLob
IkveXHUoNogKFcVqejUapHL7cdolDrwxxD8qOWEehRibDX92G/aCxzoKj7h7yNeZ7Z6P4VmBoz0O
X4mNb/vogUR8bum5fEPTkwu1BWn05+1T+80BGdw714xum1uqjF86s3cEJrdTf/RJVgwNapJzN7Ar
8o0fMkZgQB9YZZOmCoIQCHeECRPjwSi945hJZz0+YrurmD50MzrtfbMzyVVa3IZo2XHTN8G2LaPY
gJUP5YcNp5AwhsKN8AiejXVta4H4TiEuqLr+F+KRELzPHGfj+/GG34KxUYhjGKvH0OBj1Cx4eP1O
oD9ND/gfUhC/C1pi6/dyrSZsQZKwCtrxPXi67Jta33VJ1wFJ2nwqAq/IelvW19eMbBk4RIDxJjVe
WM2CliBiREIFueAPUW+8FW4ftIc1V7LjEvNskIU1VOCxyHRsC9uzucNPNVHZQgGVxoECEO/bum2C
gVE5p1+1KpszQeAlV5P1e0xagAyj6hY+7y0BYJtA9qTCDj9kUF6Bc2169F3O0x6PVpguRdti9RXs
jG381udKsE18tchlvFMbwCTt4gzvzb3Ok8f3Oq/viCXoCt0JXtSwujC++oFgQioaY7J5Zy3NtYev
L1G6Igsnv8WizIlAZZa90jhb3Wew2A06UwPDC+q4HhCe/GhqhpYxtIxl4wkTl6hCVihYan7Cpdjb
yPwLkCaJaCLsuqExrcoGga+ZDMzBTr1hRobjdY1XP9YUhrJwLd3UY9SMC9D0mWdndb1228cL/BeR
lpA5VXNrx3Ibjols5j++rHFi5WKWSqCpGt7HSRCeIzWx0FYukQZnmciti/UNd/t7UPM6rCNdIp7U
w5Pr9aeUFWp/i3wAWzOQ8qmb+2VCHqkgwLeX80s8fLEKDfuH19rryS8daPqdTZSMl82V0hMrmIsq
susv8MOBfNQ7fZl8/SC6q8z2fcnuMfSKF7opZrg4VnPupY6knvfzw0I59X2JPivIqaQmFV0M5cdT
0eR703gPm8I1IosaEgEeVW7UMlrJFkszAnlm+8BHl/3BHJirG6XlLSaYhd+CNOJ0XyukOWmpqHKg
lBAogLJK9trIzymwQ2htMkll22gytsn0f9JbpJf1b/8qO7FcN7UlL0TGBrgxBle3bF9LrDTjedmy
R1k46UQHudmWne2DE7udWXg01z5GU3wUpFF+hIqWfWiVmWV1KriS8ZEU3bGwVw0p6V4873jPBJEC
DedzKeHzSX+fRRiZjvMYEKokn+OuUKde2TdprcPknDyPFLu6JdxmjRy3FrXdfDsmVe7hXnOusrC2
CmoGWaBF+hVNdORKC1roc/LEnMqOK/OlnYRA1OiloCDcaE8PSAeD5pgl545qsPi3x+efB3FzsHCI
qqr9eOtBHejekdY1Ws3ICNnPRR9JupndZp46R+XejKn6PAPvNBqzzoBwokUNixtWl4NROQhd2lCs
GyaazMtFYR6dc5UIXv4JmEpxn6tG6OWo07F9p2w2h4BPCURm/HvXnUbDMD1QKNdeHu++lZBB9a01
cH2qqaD/1QJEsGaiVfNHLlg1c98g9szE14vaBqbKo/lmlBvxJ/IhV3WKZmvN92RqhmM9qBQkoVVp
4WioQqLKmSxDoRa0oONNrzjTcVFbUGYbH3hHDH3ZOT93UYGu0YtxWWjFlJrgej4gTiaHzAjVkPEV
VnVAxmxbUY0yvWNimcQOsOxZkHoB3LwynRNHbVvSJ/wcXC81BmN2DJRK/FKoc3Qk2eQWsgBalYBq
u4w1uZEekb8zdq/Y8cAMLDCkKEde900Mpikq6rAfy1RspoVf0oHX7X0mkhJF/lrRz/okddzc2dWY
LH7UNqatfyFkzf6SsPuG7K4bvAbdlBnseQgIPw+je3idKqWLBFP7Z237bgbiWG3DFmdMsbrBbrqo
LSxApkGrEagi8GyonTt/C/K1B3uw6KPOnPs3XcJpO1VvVXL9rQPuNgiZu15hBq+TsOITWYyThW2n
RxSwxWYWEnrfcPfT6eJ+rwpRQ/PceYS1QJ1vFEbQhpcS+1R4NAAaBEK7gZp9nZHm+4oqi4Durf2t
creO85Vgvp0u1FYejK7sbJtzYi4lBej+EFTGEusZl8LqfO+rvIcGgyO7OmKPwNfjsnJt4C6oyKGz
odtOjWyht8VPtErDOVNnF7TBdRkuUDRInvLvrOnqvxvL1BdP8y88PBbohyfqHXshUfngFmAF0Byh
UXEASjK0dDIxoAbrssi5ZIVaaBdVRlKkUCxnIvZfHVPiYJDnBut8/CV5pMlH+BzG9wfr4todjoSt
tKVHgwpu6V+7hK1JIgC91yyeUcpFefv21YrHxdIZXEEhABuC4SWoTOVtVkzNxJTTRb/4ZOHjK0MR
SH95lMPL8vQantuCz1RrD++jc28iQdDKVKF8jQfldIgscaW/XJoGy+lSH6Ehyd4ojlnrWnUOMaFP
IDpR6VDVaNB5OXRNHUcGOBhAvL0DqnGjEpoCB+VtiOySYMT6G6s/o8zLCanZ6jiE+xb8FqEeQRk2
7v1+D4EmVLMBUXaeC3e9e2fSGmn904QCKxut1Sr3OuXLR8U+/MKGwYaBqqNmVEyD/er9h+N/jwjI
4AXYn2V0A/JJ/sUajqgc7WPTSoXVAseTRR0Ce+42MyPvxt0XWAAosnt+0OX40sDqaGSpeb3u5+Do
CBSupUS3SWgCvYkd+910TLPtDH3lrgR+o2z0BZN5H5A282nDIe3Z8MNN/Uj3/ACgZ9XElf2w1ydz
EvRcto7cfP4frilDpbntiqUyGoC5Rp7uTeZzolNpPKXM+dpkzutrQ47l6P1GDWKfXixg1t2LYzXr
MaR9CPN5OL6rHN7lbfCbJRsASvektKh2n8le+1Iw/op53IHXXIiylsbxj2RPSc+ID4zqR/7FmspL
8pZHTZAu6OYs+uST1WQrvCUNkijfKilHXo3GKP64Ou/e4Tnnc9wu2R6xlOSPiQ6IzuFVEXi28mOW
iMQ8UWVtvPSadIE+ohzaIp5LEICMlVkZE9BWUrxb+2spfSCiduZP+DZ07XhjxHzqlRn/zDz1GVYd
fYEw/IRGcOQ1FhWwQtbQhzofQt/GjgaaUtYQphnufEvO/L4cXdu/udEDfOmu24ygpk3C2h6ByF9D
7VyFAnSmIZRb2g6MPDrPzhVALXWWu619c8N5K+aZnq8+2iL+rsl8nIeh+XVM+6T00t+V9ORsD4gA
Zl4iMNtmAeymJ5fm+/VA+0frfmTurJ8C5vzFFFfBPz7wKuHFeJZFDBrAV037lRUrtNbKyFGEDcF4
FsxOjDJQ4oACnYEv1M6DsDVw+CXMAi87B7Sqj8iSoH+GgkWbv0/WKsLy11L4JU9gZUlsql1LiZlh
rd9bwyU6FyNpCAosoqlXV2VZIeZyWxhiXB28eJ2EA3hZAbmNTa7+JzxsSgSi9er0S0y0BuKpH3lw
VTUeJegNdPb6yIumYp9uOeuOJjBTyfTk745Q0ecUGv4FPozYmdIN6SDT5WDxTHGAU+2+Lj4vtbQ4
NuzPYY8CNOJyitiLiEX+Zh4o5urougBJLqN2slMahTNiiccPo80qGmCMAcV4DnhXQKjXLJl24wh6
sd6oYYXcsy6r/8WY11x/IfacoTn69fJXpfq366KUNbQPPxuDhMpBB7fToqxWIP2bvyP0hnveMivv
VGwHWt6h94vr51fb9nc0LqglOBIccdNzE1Ow2H54JE7tO8WPl91zix3Y/EedIgq92w4mHb9XS+uR
DG0pS3Ii+9Ae+UxXHekzpF9X+mnWyrnqEQS7A4Wo9aCupDGYJOofAhH9A497UcGF9BnBg52cFOaK
TUGPdloTPPdY3md9tb0AAImPaTVZONmqfGsz8SIkWF3acYy/h6DHADx0sSt0gtqgMFfNwvGNKaxD
lBQ+aw1YO7fn89+ayh272ynfsBdOcpUz7jYdT7SCGnYyDOS+V0prV6DyW1H1KKDxY55YrT8KTcai
0tJLwXWLlZ5oVqQHkbnU+WCeRD8Aruep7s6Un3Seb0U41haLm2XOJK/yzA2zGia54v47uZqnWOIe
JaV8qRF4BIbtDkNgkzpjzW42FryGMB7DkKSultr2rFhYqYPmHatH11DnNkYyfyQQEhufQPXTV25y
teBlncP0O0CHt2NjI1ZzXRRrEirJ17rhxk8/2ITW3zC62bfFLYChIxLn+OF5cg8fviD/uhl6w6Ve
iaIT71gAMmZ8UUZvGKZsi2Oxs8/a3CKr3pSIjljz0T6ggTrHyCDphkKVf14+xQXNW8Hkip+YEiRg
A8iy2scvaJIuqngHoS0RDrjB1ge8jm8NfaAnkrFJiYm0dCSRd3Goo2cp+Nd5ghsFj2nskTDjt5hh
h5FKfyPcfX+7XDEpmgPYyqQqBQ7fYm6k/7BbLFTk/mjwhbYpMMgrZp4OFCLvkOy3j1Vds3y3Cwzz
XV0HTV8LboXB94rruNtuhb4yc9fEY/PpUB9us/3E+AYRqv4kpe5QwsWZnUH00RtsAGjTAnwEqfTH
y3yM54MIWAVl4iaKRxSX5GMT+OQiLIRFV/wo/5qp2MCmEl1DEpW04Pob1nEEaEN25VPY7H5xsHEU
zKASyv6ywDhKaTRiGaMsbloTsMHoCc05Nv+NNQCQIN9NJadwnIApzNps8NdR16AiMGPsYneWfuyv
rpS6Wk/iiiJsuJQVz5tE/0wgyF1onfm5tK+bdWhhD5ebRylaQK4oXE+NVBEpthRRoQn1lXmZx7AO
e3LlSnvCC1L4os7Md2BhF7hJc/RPIpp1ieiUS6E7gE9yaGqfCj4S2/aGQQ6t9jDFIlrDqHBb5BnA
hPRT31LzDE3r8I6t5IQO7MIno0S7huZlzgo2wXUntjxNv78kXHpsVGG23/vmSKbfMvm7UQs/oXi5
N+XLE5p3mxrBuDekIBE8+OsdquqYuAOkPDw+uWXDHuLOWg5x8B74pmUIPqMXT5+gfhWZOiNrm/AH
DXLvM/KUx9d083Gsd+5vjxas8Wl99u8FDOqP/3TkU+ibRO6w//Vk6xvs88cQavGg2ukzVlqL0REE
aSRwES+NZ5WIHv1r50GoTDwvjmQferJeucwfGZJbg+/moRxR1RvrSCFp2+eSY+7pX1cQ4tDQggcl
nCVfn76Mf7R0TjSf4rYgoGirMynQl7Jx+cFt6sO7GJIqh41JipH1G0GMGC7IBBU7M/F/N8hNEo+a
P1hGIeANb/HrMlj7aH8F3UVsz7vVrSw6dqB6G8wbuCbee9k91YRLQeaJDuOnKwdw95/UjHxiBw6t
DOyfflaTboVUiRYdAMbWd2huY6xKr8USERyGnupzNeK9lix/ragq28g9W7u1KuYUVwWNlM/h2ymR
wPLfU1mDX4fMyWyuTbeuCO6+orc12ZyJCgohrCQXn3MQdLQxPw+9HNgIFNQD8EXPHWapfysN/wwM
VvcDl3RIOSP0GESbcvr2hr97sbJyoViue4WOLiqt8Mr2/GBemQjVMrSl9UccMEjK/Z5aniAm3WS4
nvwwrQYKfT1J3PK9rHWrVcqh5Zi6nWDJD5QcOW52VUusA/qn9QMUSJLoXvzhoK3PJVzp9kpT8tgn
UWopkRKsp+No0qQQ8d1+/Py3/LFnG2bijr4QQIN4uo9nJXOV+zItA8jriUE21///646mmtUJE2Ox
U7y++5yrUbaWtthNE5BSlQn1vO7fUyVO0wdVFSGhNgxhhOahLgODoWF3iEfNW0jCw3dIpbqkkc0k
uJCWWOjdr6wbJ0oFQ7nGPEpG0G6vG6LgzE/HupBin6MItfvG1763vBNds1ih+KGmA1V/lOwB2bmp
TtMNHcXyxB2BrFvr0cFp/dtABUCs7+JXX/m9dsjpd1+so1VP06jFdZLk88T3+v2vuWQag+M0h1S0
1A0BsjLtfsNReDEy7V/qUDcs9McxH4r8Lucwe0+OsO6L31X46hOfKOvz2RY5RVj+rkLrC/pjqvU9
j2drsXm9Nye8kgVlDHTXd+GK6JMB/Zv2FfuC2vs8wuS7QhI2eOc5XGyCxbGzXcjoeh/pgi1JpWw/
Ik/CxjsoooMqFM2Ehn6DmtGxSpltew8hbAnWkR6EyUqhkijiF6iws58H0NaBPaU6NNH2bHotHQbP
HHvMoIHHYPAcWPKpCS4u2DdgPZmjI1I0BDNodXD1ALlLf+I57xc/MMOv+Xao0Eihl9+VhQYV5A0M
R6K/6Kny6ACTHCXkxUfeQgC4P9jkbkb73bXAHjeDi9IprTSTg7EY9mNGlwvI2k5/u6C0moW9KvcO
CJfu1Kh1zdmeUwqob5b0Zv/2ZCEN2UAAkJG9ffa/G+o+nXHuMTpzXH+RAPhMzH266S0E/JA0MSgB
wxfB8Lz1kCDjNEthxDrWYCh2B6hEDALVgaGQ9BrMwFZgaYXXt7svyb/hxQkMjY0Qmba/DR6RLvUt
tyVja1A4iv0KwMprhyoyHGP64xcfQOZvbGuJqcVJbajOp2HnfgmVVX0Vo7X1yaZzh4iu66FSZdjN
XsjSKr446ptENohF966+Jlkq4QG+QuBDEVHuz84PnfOl5HEqJ/TU6NA83tM+ttVoOu9aoAv29+VN
Zxbwbuv2LSETba41wFsK6CQminDnZC/qJn+9kVEsRv9IgYVYfRBO4pl2tCd9G0sLZkHcq2Ll2d+t
tcyS/s+YoiCZMD09JVGvamF+Ua+KnKITt4TTIou0ZG5tTdyEIE6jOJmYc7knmL0mFk5bkJfk+5+K
O6WrfQfmtvZcGmCNbtjOpSXCQqLWM7Z3KaQtrcm9FdC/IeQEzHK3m80m9MI5GTsPW/Id73n1GRUM
xg6j5ZyhYHGKzZc00qlSwvdqZOOW2HL6GaGNeB/teTtfkUNmHkpHBqFnUUEtxwupYVtH9Wn6XjdQ
7qTZC9nHqLnWHh4iEl46uOZ6l6x303oHJavOCijCT0G4LdgCIP+zcGmfnhgMTtfYv1k138aw0ytb
BUPFjpDbgAMoIatJHkglShJe6iCd3xoO10BlqPiv6Jszvz3UFkrVF8AN1BiZX5jClAomUvjH6lKt
wm/yErrLZyPFwhcaup966G0sr7/n72NM1vBOFKmVhTiBwR2FWOHk1dOcPbxvHX0LvPY0f7HcRay6
PCWSefJ17oMxdkP5WDs7PsGLKxcyoPLYMeXvTggeTQZxikYRIu8Ml5QS5gCyKWJ9egpTPgsuN1vV
anPpr+jNx4u/08CapBgz1I1GW2ughPovwJLXruL2t/nCx4RVLibrSpUaksl9KzlcVSMyUTKOuJUh
D4bqx9kJ1hm4z0IE+qnJrbSMIj81+I8puZG2KfnNz+NO4r9daUd7nFKmEH0Gpd1rRvo/3CUrxFNw
h9y0uO1zZ95IEEt5VKTou1PKqoHKzDhlybO8UkbM66EZpk5/BD3+f51499fYKI2WL2HFlHrd17sU
CaF01SN5Sbgg6djjJ621h41RlZ/8w0oy0ERSbaUUaz7UvqF3SR3c3GmEJAxmMPZ26L0qVjGiQpxw
Do6HVuUZFCW9ptDmRt95QQjp94eJCfZldWQdJFHTg7cnp3QZxbWkoJ4UaPaJhTebj8cRJbyyoASH
RY2PcZaxmRwagUiWsWY/pdd0OKnnp/n1KKqTYz4wutRtZ5+oBFh8/EBJ+mTh9vv+HduhPI95DRfa
CE1x7s2WG8V9SOOociw4P6DZ1qL64zwnJE132Ik/fKq0Cy8rANpG0k2HV8gEWeG3ylzEGBiBaFji
8P0SfysIGzR9xSz/HrErp8zktD5hkBlg1pwXBqKGKdKBHv7S2FUEak7Fm6taRm0MVH2Bqa0yxdQT
rAvPsxlrR9l5Zw8xr8XTAzodTg01AB9IkglhzbnoHrNaZ/nFNv94b6qjZBkXDxgbnnXTBvDTxQAv
RwuoW/4HxQqMzkcVtTQ00puftGdWh9pysZs6XXYNYQYm8/kK+7rF4gW95TAcuHYl9+C53KQeLmxb
LLWpy1qCF8JPsjeUYnO9FgENX1Oss5I9eZSi5RsZCZiQAe5aflm/YBPgg4y1zLUN1vaa/XH4k2PI
XIBDhwl+xz66GRIxl9YPRRS5Qfb6n2JHYTAwdGIFicfRrlW3UVXEzK9yXx0iaW+IACbPGNOSF+pV
4jGmDBsa/2K99UJYR49IgsecER1epXheI24UwK2zzntr0A1DzaCOWZspfwwkAEGYALhFvy/a/cHS
BAbIxwBEr223SfKWO7TQ8UqArYG0xLqbsNc3L3kqgIOF9noxAwSPPJOFx7SMDeacQb2OuK8bJEae
FUUgxkf0xX/qkaljXe7vVGvDZkRbwM2EB7VwVUlstf4I3EuxCGKNLi++ghUNsK6xWeftu3AixAqn
MPNLQASfk13P/dPmgEqdvDU1lKT5Criy+0nWW64mw0iB3v/dJynZd6FymjdUZv+cGjbNvTBwd9HY
/f+kqayCYOASEECDqPyjydAUJDGy7xDqhi6F+bMLkczetgUONjnDzmIfoqoN/uMnbhxzguhV36a9
if2k8M8L0dxmQ7eFrXYcwFnXv6GPx5m2HKZftbWPgr+2FYA6mDXkcThztodtMojdxDvkhLBrhMw9
YU7tPDqVJrGcq8KPivw2aR4qo7k1BxQsyH6EosH2k8LqKtfSutBIOwcqt3I9eZQI8JWoR5w6XCzk
j0bWgsYdoedwyxsLh5+IWawEPlekuFGOsIfV34gbSEII+2uVpZXRrrvLk2w4AeqQ/L9RbaKmiWeU
ULrUR8syIgeAu66YTBh9JtFIIgkorJPUXg247pVPFZNx2i+Nr3wHGYsrgRQJKKvqkaax80wzpvw9
ZtG0jy0mZMSpgg/3v6WJrQ4ulyjuMXcOmIIhYOKyHv7NFvv4v0+WTLibjxrsNEvGrqY6+L3+qX29
6/Kf+cBCcduVSs/MOKIkFhd4OtuZr+6K3IZyPWFHpciGj7vW3s38eH8FbXva7oqJ+Y8PmX1H767i
Zk69hJhwOwelZB1owZjJPgYqVxZCmUNClZ4Tk89mxEnOTdvRLwIjSdLylqS5Xr4xwVZ7YQ3JleY5
so/dUAJ59IWGgBJaYzeySTzli77qOtLTvusuGCWxmia8wBdVNxZ83g0qssYZls24oKbUorSZlZaV
dqKiYL2t5tWF5MjffSGbzSL08Xem2EUfpBPeEDbt/ti2Kbs3nDB2r7HSzO7vHGlouJPHR2PwrQp2
37flCl2I7zObATZ/QL3/kVjMEVOUdYLBx9LJBCY1pnzRujo6tjziNTSz3FHDq7ya9JO8Dr10rkrd
iVb4ikH3Rylup6be67pYtlAV+RXzPUYQjg6SRttXTWVzyw4465+FNFhtrh8VtljRz+5u2s1He+Uj
5TEwht0bRzvEc4o/2EonVWkYf2rDIu1m3xJa5zD558OwvIn0E2sefcYTaq5DEhZzNS6bwFH8BWc+
CWIwJOp+nIQm8BCuhjH/m4GNrS05qyZluuvseU14APIXUWFoclRraP+9fZDhTU/ihAe6PCFCtOLS
lOygH0UXVpr517sum3aJiBqAL/zFLjtrtKqWq9nOtR9NTC51yH+/7LHhFRyrDPhHNtNtnUe7kboN
6LQZ57NzxSicPz7trAomnFnOTmnD4cD17HiMFCeWJ5a+p/KyDAWPLdl1bMxDo4WpEktAV07Vezot
UnhtPnwsmehk6W/5oGlwh/YledV56FZEO4FBIprCiEgDOLijkk1Ye1S/BaPSNAnbpw/66iII5CAl
nk4a8f3iTxv92fXjuVzdgWvOLBqf/c85X2e2Q0Ywu5nGr37bvNWhJg2UjTRZI82iTepRueEUVwCO
gL0X3ZtMLzVCoEjVCpK0We1hxZTx62ftEIoCGuj004elEKuJjOQhkKDdwzz22nvgmXcZxIE9p2iq
CPbW26ROuIHmZR8vSwGHZ6COuejkSpOr+SNjv+SlDu4/PwNLfSSpUenQ7Rb4v5Z8VQ1xjijhc8sd
6M0hguJKZdmkdR9pryjsvxG+6vLYppz5VQVs6wGEhmqyD+iWLCZlTRWK35DtT0BiLflHfsSrVqvi
7+Qkne7LIboUFav9Il3bhBWDMtyqfuewzp4z3GxYoeI01x0F/oTW1J4iHqpEoM64Y8vili90CNXK
9V2V7DDaagiup3PWgCqR0dUOoMt1QiLVBtD4bU7ud+FLrEnk5YQStjM2AEPMvQ5QwW95N86lpNB+
vwwEXs3b6uFMyyyNUCD1FrvixESSf5ZXzEVigyhHNZ8h/pH86bHNtkvvcom+1/LNMRDhQYVnpdc4
jL+TW6coyZVOmo6bUKjV1qQe6lklahUhgdTPmqy2WP4BqyNyWnVOlSnEo5LjTIiwfx7tYd7f0TgV
+j8dBE+sxalQ7bJcQOJusTIsnK7NXYfkx6qqzdYruCNqCmUlHb570FYRRFBicMbcqUbK+lY1RUnz
Y3c1Q8pWFyY7+MA4HILUyRuVOeCiXq7TrzH8EfUF+3VKdv1S6N2fOKsOfL2gLid41Y0ukS+eH2mz
xrClGJVPPKNnSS+NlFkI2uqJ2HNvj35+pyUvUe+cl7WFSFuLDtSIR1Sb9ND6WNXJaJIKCcgDbceG
5L6RMbPXcdmniFnyfnFnExhMXB2dqWBlvLnKje4rYeIIPt53xNZI8hwJ8f6oyhabvN1g25OVMIGh
ye21hz/kjGKs+AMwXDW9Ct5fbhIwb0nSzooQgdspdga6RAiUReNFUsMnOn1BFrYH4kx6HiGUmzay
drUT8SI3emcqzTr/5U3V4F82as1mi7593lC9nwssPYv3mpa/klrkfq3YzJgF64df4qjC4G2N5cL+
uslDEcL9A9/SWNRtuNHsm3DeDzXf+9jxFCMOuCfXBe85svwpke2f7roJere0RcvjArbtLvOV2qcK
YufFlZ8MqgQKMKagp5wMv+M5bjUK2zwq/F/4SrLPo+THHAzXDZ6xtaBMbaZSl/h30ZS0ifiTRDET
+CUBeQhJaNy49ipOp2iB0rSdqe6mmVymxbA+MFAtykSXLnC/SRm2sdDBrBiZBM5tkqLBp1N8kNWN
lsRlyqm+2fSppQ4uvEvHIhRHbh0XFpBGtU5sbx9QJoOSauUPC7JvOvGPKHt9FpPi2ritEXDuzXrv
YGG893ugMs5PcA3wiDAJaq9rBAAAb4dRe7evyRIWtqpJT3Ng9RwshbZyGRLLUMLmdNUwm5wUgpcn
BdsjC9xGC3K1qTTe5er68oupVCSi4sueF/XaD+Y8jb8rq/OYKaXCtStM2UTBJBdKEacc1FskPfgz
hRmJJle/21USW3aJqotD5JYIRCAHd3xk+iJob42I1+RuwYvHz2P8ckhMEZqVTYvUZXOD/nDb4G1m
1TPDqVhopdiTQ+6+OWN7bDD1OZ6G8w1stzamLfEAQik/7+YCGvtDVdcXc4d+WvQVJSgnNIMACKh+
tZH6mtfNVRhLara1ZB8ejB6PwqWvNKA9c75yxDBMQJIV1KkYRRf3ylpdd+Hkz9GM1ABtGxkwng+R
9VfBujedvcFU4PPgXHLHmVenv4HBbhbiO3tIjNy8oHp/HBsMcdaCbW5xvm2zt7Sddwvgu3RHVVKZ
aT/eZxMYTlq5MMbfkAbGjYOqf44HZvVWSW2r6+qf92e2u0t85MOA7gHwk4DVlxkAQZ1VrI9aGW79
MIZaO9CgqZXmYbDsWlqTcjb58qwHgnheH/gDF7tfCPq5tB9J7L8fLly7z5YW6yr1zPJa2j6O+TNq
D7phUrzTSpWvKrou7KXD/3bS4XS0oqSIjr2OLNnQqfUgzLdpGIVRT+YiUhaCj6cYSX/5wqKNV1OX
8f6IZNWmARld8yy1eETefdVAxPPq4gqHfHDbAU06jz/ra1a24+4C0Jo3JTZ3nN1z7mV0lOYOFwWc
DvjYScm8/NJKC1n5ZTvSPLAiF+oR0ufAE44d5fp6O1jNKOTLyL79Jc0XaIlVzlZe/LqmA4VwGA/R
jr7ZN0dIxu76R+7X7Tdlnos9l+Qz2JZGyKj2V74uKjOzOMx+b+3JqNs08uTgonXgB+gjDCc6kTyE
Ca04+lt7uGYXqfx//6KZc8GzBvB6vQbGgwIqszn9iydBTPPkTYeegQ9rqXhROSiXwVjJDTHXRHkC
ZoWUD1jH80qBBgguT0SaTq3w3MuWW5tlE/4Fg42DkUv24iD1N+D0dGzduhTaNjctEneawXoZXfO0
KizcSjK0+h9EPohTtJGnv9P55RwBNjUfMFl0uEVjxL54dJRqfeJ0gdu281sj2yyk6rRJJe8bsFX9
NlEf29e0pJ4qiV6zDQ2rWbM81d0xCX4XQbpcOl1BOdhk8Y7MAHPa6SQywsybwSDGgBSkpDtg4DDH
hvF5g98nvRQpmu2490K/abmgCnyLMx4Sm12f5d6q3lYa+EKIVXWXew5+HVD8YsRezvGTWHjSczIP
LWpCKZ7sdT8yd7xwEQeH4WZQRUYCs2uuRENXuThMGpgG7dcjXfNnYC0lkx14ZMqHT5F7ibZC0Q5g
rNP7bffbIoZwhZG/aioBzEnogxqg+q4FJ4/4grJkdABDLB9mrwwA9CyXu5t7Wpaeqj36pVGw+Um4
dB17Agokmn6KOwQSKOgaACaefrfGg9Koyd/kR+T7E/CLZLCJor9hH0jLeQYFv7jVpsTBoz55Mkgy
tytsPB3xr2yUW7+4xTUKEYnDK45J1IMrJ/PAsM+FR5sjUhTqkAzM82Ct/cHnYxL2ekpidR3C5IN3
wxYWzra5SFBDFgJxmWSrdro3xDk/vhTt/ilBBtlwUtbvftwLBKLQvZX4vvmTan3hCCF9e/znOA7e
5duzvXGhfgUrXJanX1ThHZXU9JxLAJWGrySQpOG9R8/X4BNUKSMnOFVMrymae8rysAVlfwlthZmx
S3sI87z7KkT4M+RQ4XoFaRkdviekgrjIMxTrkGN8zJ6MhMTE1z+v2Pnriqr3qxbUSiRELKg3OZ10
qZluWYuWqGcgq1FfPyCydEK10pFh4t0l87nsPgwkRUr2PuNQ5v72ZDmWKEloovqt9uJzeeuBnoUp
/0a4Hz9xrsXzFPUn6JybG5eebu+loxp7Uw/eCIQixTcoLAtWiaaJ029aHaZs2rKJQxLNX3mtYvjn
SyRVbTIF8I1H8YWKPy0SVP/S0KWeaBCIiAdFWTRzXtknrOVGVcQtmFWhrHhBbxnJrEDc9SHAPUAF
989LxBCYVimdoAUqOoaJLaNZSeoSBXh+fSxjr7XzICqWJ1+dZI1NhA4P3K8rLafIMlAuywjCN7wh
c/KDpy6tf9AipqMoa0bdX0Ws51H7ROlnJvaQ6w8LkH/AvNNGjm6+iwXlgZF2O3hKaNTkw+Gob4sB
lCSB4zdWfIQ+jPza0xSCN3hZLCsQNToEpB/YkrWS8/2RD/GLUKpoXjzS5BOzd5q0ZPIhjqeXkI6R
C1H1kefnFxMhmBYFefEHstg7F4H3cJItMahaoTTyjQcABlQthJrIXDIDMj/+3CAw4B4Cy99tYwj6
Xprq403o2JDWWTh5YEdSyLAjeGrdfCi0LV9FzyPoZq38E9Or+NwC113eRkHArm9BvR92//JKKj3O
Vdxybx8ErpTY76nvgDjHPPql7FIPXUFXu33PIDzxHo9ymBlDmabmq6eHrWi0MKfrk6cDSgVrjrxO
Ci4XPiE9V+bwe4c9UFc1xIP150C6KCYqxWkCeLfNgFzGzriSiOt7tK5WW5BJuf7RqrWYWLP1IFPH
LoP2QkPVfiM4/Uu0mZmPNJ60b53Fu1BhZZfDGXxvhh27pbzIuuwbfJSCBUJqsPSQSvRtyI6/PFQI
tR/8p8i0yXOCSHgBp/krZtrAc1EPXMU4Cvf3zytPUv4FfeL8GogMkZ3hsd+2KP9G2Gr1Zq0dYRej
QMtJNHCDdPOpyejt/q8pKGthq/qpjUV8UzdxL5D2Eq+6yBC0VkUrrAkXZ6ojzXVFIqSFdIRtbF5a
4kbR6+1WfkuKLTwBi4pCZ2JD4hDPLcPWRHGsJIBF6ZDOEqxDK+oUKDKX498zQUbuVucthNJLtYO/
81snCxTxnDEX/ImvRfEi0DplWy+/oy4N0vCNDgvY0xf/t2khz1jK46ouf8dD7CY7SliGCiUByqbx
skVAuIsG2Y+QjLQZTaHHlFTyq1O76VdS0SLcGoQq9JdLh09o/yl822iqcOlcnOUPhsdD4vz8G/dp
WFKluoTIWlQAosWJCd1KLhrU2HeMVjvoYHSnySU2M+KK+Q5DjLwkM/bJ3kIs5kdWO/TRWx4NUT3v
DQDCrvZtNl8rdcrCqpjW/7/1FZhojj4bbxzCntEBG1thLnzVW4yV9XOctGZvK4WuQDlBSQsopQDm
eFnSqqbh2tJ7VfdAl5hlu5R41pW6y2VQRabu+Tr/KDO/dy/WncYOPca+8RbOfb6a5aLgcPe4uLo8
pr4JTAKl+IwgLt7CpeioRDjYroTA4VwV6qTSActJVj+2ZiibodVeR7S31BYHL4PobJbDVsL+ey3A
nwh6eRju2MOkjryDsL6vr9r8T4bKUsyLil/euRvdGplWWBaNOGclFFxk/pJ9no69Xx0Wou78xg3t
3v+krVE9S6vJnYLsMrzcJXPwhEEbEMJl9lBbP3geIPVQV8HAqFYZSfDFSZdXoD8ZdTDpIQRwAxWk
WZNU+nFP7uI8e6zbobPsS8NNwYSUV4t4pNObVfLEp9WyOPJ7ubb3LAyX0tw0YOiPPWHSIe1pWyTB
k5rMPQGlFJwCULYvbLcW0ubuaGsFz8imyxuB+4ILGBpxuECTQfp3evM+vElu1wkWLM6kNazgX8jg
3iB7GP9xbgE04mu7jV8imGMYHFFzNCFk8LlLNtLvLMb40rQxDCE06ENxL0Chx9N8RihvxtQS3kLM
+gH7d5aeExmQzt45tKh4biRMdL62VUkGtA2L/S80//1cIVVeNQaKKqc+Bkckm8lZJH7Hvfuxx+co
UgQaONrfsf8py29GLn6xBKPDpX2C9TShP4IJHn5IVFJBjsPOl/gmx6e9EbyzEw1krVosmUNf8J0m
/YjxsRK1IQxTGdEwd0ulXDrxUvBlEbzv8QMP07ZrKUOf9umGY/opS5Zj0vmbNGTziaJyAF/g07cy
Dve0EfryOBV7EzCK69KJfD5xdEkQeKpnluIjt0y8dlz1gkX4XKRZh0iqSsizYRqSkqVgZ9sCQddd
M5h+i/22Yao34trGmCPlMv2fOx1wHPFT05NSGdZ2Grdlj2Hz6e1pvU+TT6gghu+ZBZZSuxxpAQH4
akp31CCl0yvMbvo9ddX1VVSB4Lego8YyUXf7cN5k70mC3PhWGXGdstXogC2iJCefSjbkaqq38Uzd
R2eNrgpMk60VAkX78mcuSZVpl8ctVaoiFBHVa72DVBZdTuMiqYz7V6eMlvvBI/yLpFWFBVO14HGZ
Cd9G0vTmyH4u+j4K80AvkNZwM2sj5LglBAQZied6LRgNnNHisBAymkvHDr5pWanWWkKmocuTzIlb
kId+2bTXvdNds0CQek/f9v7pN6xt/1V0bFMNmnsJmxoIHVz8z3Un7p935ybOcmrOHgD6m76rXrtb
7AyD7qUGzdMekYuG4Lm5QpgSiSiYu+RJ059HHQbYf2MWM2aUn3TX9lGlCKOAkhsUUR5/FL3oHPC7
mu7wvt/QmmvIDaIzqNrMlEDg/cMO319SzJWGjuoMBwt9//yNHG9PtqW0LrC25vBBEzZuv4HBt9wL
qmZf9/uEhU3xu8xnH2aO1HXceExNFxdRUjOVhOaIvApJYQJiWNrF1kxvfboM1dhpOtMA9QWAECBw
4pltYlsEdi8BT3Xgt8Pqn2GbSu0p+UxAbD2C7ViTPvTQcgz4h3CMIYcGVSLpxzqWOGyxbaGsWK1S
m61yRpNC5IHAPOXEbTBQn3w7Yr16zFl9Pgo2GfRxwV8rnnVfclXj8IItAARPfmAyVFu6vNWMPdMV
WU1Qr7nNA1LFpjwnVVdb2posRAcQaWpPEquSD0Vs9R08vsq5HsYHwPclibEbPn0RasEBzITLXeek
05cmhfU4a8BwzHFvyvnIp0Jn+JwOIGVP8p3hBDS5AlBr1IsY+PAFBfEJCVrzOLKrT7jW5gIdLdF8
g+ld0H4pJVtyMK6uyNX4WmgqDsxWOBVX92869wLLPWIIuwaZSXPaV4WCNv7Dq3gWmcaFeL8e2cQz
3/8MfIg3DY87MIp/E3KrBxx0B5aqsxDfr/AkMHZ3NX2QBZxutP3NLOfcf/MSCiyx0TgZkKNMbMaI
5mwOdXK5uvx39MlHKeQdP9YMd4YGVHvP/n5Jr9z71xyxNM2b2bL9aJlPTJ3FtpJLHnav6XnyiJQ3
1jgYQyZh3I9DJ06HauOSPVSRh1ymUJ19O1pO9hTnntZXIq+AU7dbL8we6idXKRhgCWqEeeVinIK2
HxWont8D2NfO/3RDYdktAl3rUWX8zPmdsTn7spAzC2yxK0NfnDZIsi4Fm94PkWG44Sx+LcvA7E6h
Pw8N9d7Da4czaESfSyhfzVmusSgM6jyKcVizRCOxvBHZMF5JamZ3j/yBWrKPCgOoZsX7J3kNe64Q
nOAAkyTM44zrqA/rTqw+9H8T9MZgHqhTgYtTpdL7HdfwoHwSIM4kUa//8NSvEwX92xZnM7hbGo2+
gwYk1hNAmnG/2VamBIZiy5RthcnPHKUx7MXzrTdqXcz0TVJLfzi7kjqMTHfmtsldnFiyjAgb0sCG
6QDfkH1FdKj8ezp4LYDd2eMdiYCtv5McxrdCMdDx4MrrdmJnyjSXG6EyDy/h99Upgq+5iptdXMHW
H4bsI2v+N/oe0sMr1rMW0APLc+X3jHhJoJLjWGqRb5kIEN5MPPDk50YANVMjsXREjjIPLRGc5PRR
rrXzZ7aL1mLLxPwpZc6973PH/b2xohgaLX4GM6nPsS7+6qK/jOzRR5mZQ0/W0LIsRK1FjsAajPv0
9VwS3HaNPLrTmfzgPEQjBmF6GEv/FkaX2cXbNR9PrR1t92pkM6cCenON9JWa53mBAesrIRIzmj4p
9VPKC+jVowjiENhv3ZHq6blfEh2p8AaEp+099ed8sGdM1XZMDwFZGb15PJgst5Alu1TLPEZD1T29
G38ryRsAQ1mzRPZX0PQJkGMOIAk2RW25Dq8OxuwTHiq71oH3a92uQY17hN+QqwpokbOqp95S8hHQ
h12BkZPi2rngXn5vvb4wlc4HOjRXCrEE3TmZZPNVuu3dU/vTti7RIq21+P4PTZFzkRC48fbyJ7mH
HtvujC7LM3cHpJ5Qe6Vf1HpgtnjlgUu/mShAqZ8IH6bDdy0UT8NzHUaT4gMxWuWIi1R2amvId46l
sKcfdCTmmkbz3eWEc3046Z8cS7g+zFzXCBezFj9g7RdTqUgqad84b8R58Bh+c9VPtpaMspMN1DFe
+G5D0Jk40uZ4HatuXtFQhlfY/fJoCDpqFBkzsptm9PQrmNoNKXRVaOcbr2JaCKIvHx+GjAvTs9yf
r6DV9oIa7SEo2qfpk+o7Iz6l/2Okj3A5BCPwHqDw2FI1NXn5xoxMnk6EIcIdRRPI7MjPz88MmDbg
zrrhrSKG+PUM3Gk7/fhBeFA499WYSdW83ek2OodXS5nsu21KQUWJ3ozU3MQJsPjR9bXxDixHctcc
66m+iMOD4eIT0YCGLYrYhT0iT0zKAEGdM1tVDKLnMkOoOgtnDXJXGpci0qwNV1xSZG+A/R/PQDVK
MmLvtzhj0DuinkPTilunXth4O+pBgxGOJM8i1EoVmIy387IC7ig/u0u7ugx8icRz9z0fB5bcl0YG
PfOHDqs2AxHLsnL5LTxx7d/xUc1fArNL6dGzFPiUh9qMZOoHG4bRcAU8zkcqZLD1nsEPLshZZ3BL
A+0MLOA07ds4mASJ3tg3dyW9qniWd2ThoJ1HXT1I9DXpD18yapLb8Hzl5cO7dzGQmVK8z2ALElpO
54ZC3/BeHWXug+rJg1mCYYezndikjSgpcFCVEzLs1A06pZdC/afp1qTpph4nGorCekVgiUY5zNox
ydZifXS11YV7rDUzbtEp1nBe1P78003BrzTTQeqOYkvMoeXnJDDJSlqg+Clm+5nTuMQtjTUAgxRR
bfcbmiN8oWoumTAIkFXAgwKUQTpTOVgzFOWahi2QQZRCK0FCw0dd89vpdcHkNrgwaxSXcC1GR7v8
7fhq7ydmIKUC2/YfRncCTMhl6Yr/+BLZV3TpduukYlsrLhVVFnb+5dTb/ykweH8F7/UBwJMVEjgE
QbjqT+rRjHphb7b6vCqPUFL8bMI+HCEAtxP4EmkcTzywdt8vu2mmED7e+ATzL4FmxODrCaQslksM
GvE/naNdGi/WqubWBq8g5IJqjk1/fCiEcnDpnAiZ4ug6hYmennpwvBkXj/o1isfnpgCCNAQlbCha
3pXRCpm67oT1XFL7P5OOqQ1yC29aVxL/YCYN0g0uPSibOXW25EfDUaSCM1Sa1J7d7nH98At5CYkE
lZeWfIKeubhR2Q1Kpcahb+BDBhZqi1CmKTTohxz1RbC2X3f/l6Szy7aut65yIXJBhiJsZHVxvYou
bGAjZFzjN10Xy36Ot7xULivKGi28Eu6QwNqgM3DYZyX8qInKA85r8dQMF8h+jXIM50JKpKzw5gfr
YzWUpQrf9LjdQLkM6N2I5+NfsF9v+BSzNCvVuWtLmhdB01WAcoVrm+yAOyW3Hd5XvnImNnNNZeEk
JvBtPuUVhJgArxq+M0nO16tuN2DQvQGra2UyNDNnef1oZLjBN3IcQe62zsViD6NFqqqi9db2nTjz
wCMCa0nBzansS2U7EarqIRwHAAizYzanav5LWvGekIPDsVM0vgWlxVxa8EHg4UsHhpcmpsi1eg6r
LR7qQDIh7pdxbf67GWqj2pBtWlX2uJYsL86zIds+Fff86N9d+dAdhDk/nSEOxayRsde2NVpEQ7Yc
iXz/KEghzlZjRrqJJJoH3R2IEMijJUDXi6WSiBA2uhLNsibuxqw1mPZZiPznKEF0mzjW7FVvakB0
pj/rQa0a5GPcI30hdFUH/yfEyYZKV8MSKcoJrVVafl0aKaoNq6SuvXCQunh7dozIbMrw870zSioK
jyKyH0ULVGML+7Rndu4M9knbutdpuX/xF3DcZoSy4zGHDjLaCINqM1guMwGhQS+k3cOiT55qXoJY
xtnGO6vDQzFHA5GQ6m53gWyGznx+kzSEVtB4F7u6aF+bd4VPOMivmGEi6moyQReGbrkqbmJFvssb
gIypye+zXcpts2q7sv8HD5XISplqj9e5ftL95BFbvOUuQQfsQ5gAQ+wQvdDppejtxrs/EW5zpwa6
LSdFBO+UZ+3HcvNFSjrjstsY0KwLQs43uo6whP/siBzz2E5OM1MYTb26vDmj9iaHYYQubgW3sfWM
FYfgcAK+MTAl8rTibgi6JvuTxGBXWWF9rC1DFX2wBmvJKWHV3Ks9MOiWEEL0raEJlhJMAkKLcVVD
16XKyHxMWGqDnjXUYYrUFnP2FF3IxcUMVis1Qyhi3wX8H59ikdEvozxJp9detEn2PDt7HEUHOXvV
IO+2oi572mwqhOECL6Uo+i7TfuGshwGLTmhpCqlRQd7xYVhH4a0pFOSmjPmTaFPEnOhLvtxy+7Hb
on7Ako5qsQHhaBpjU4tIg8eijboJh0eR/CyxqfXQa2np7SYbHogRKn6B+JIQgZvoyrIq9oPYZHaF
KhH9/oqhDC003/0UgoYqfb7cWgaGC7g/d9PIAYYGdjymhQQn+OV5odaApBQopvJhJI13XReg7V1q
mgj+wtH9nTmsQZfp3zP8d7JLuSP6p69CF2/Hn7NvmOtFChvFnxZFZx+9o3Wa/Zjwk0aJM/T6iD8W
O+DbWhyT5lA6OQ1tbQNVjj7MjxGTvm/6Xg8G0zu3nLjvB1V0xSb4dpRQISuS/BgEFGY+XVl0IHBV
YahGMYUy+Fyws48qlGIrn+wkpJvqDg1ouuwksELGBBlyT4++wu9FzD2+rfiCWeUH2Vqm/lXksXYi
61Ks5yMn+x1ca51KZ86ctTpahToQuiAnAy6dQdKACMhEkfpVr5jsK7F3w9qbm+uZjPQQzDsi0Aih
JPOMo0xDOspSbvCZjktcl3bf3hT+VDzjvmKLxhKWnpOIY8tAS8Fl5pu9b5uHEIWdl51qjbK6r+zE
ypAT1ibe5PkE43+9l8gmfPftabJ1Bq5T+nuLkQLtwl+V0SJKU+w47E0swsbjhkz1NG4ylDxBwPZe
pXLWoBVLVZY4o7sH1xl9RMrKTPZr9JkxT9sSm8fDalSssUMJKgtLsI3D7zYIBfDJ7BXcaiLjXGit
p1jLdh+jG6tBcYoKYwaFdlwjj2Sp3ha+xtj2PVR50t4EHKwtwrrtmcnJmsrsISh27l166YxB3CIc
U4WjHeIWGFAxNnVg+ehnIW6yTWPkB6hnHRbBQQ4o4mffaR8HBi5T/sVr14zNPCDn+DRxrrseYgT/
j+k5x9n73nnhFzzrx3Abo+AJ3wqhgEYk8ZXhkE1uB7Un8Sk1KBP+hWzYQuFSZEt1A+Ck06DWBJT9
XQEvK+w1TVHpNrmpDXlAaSlkx3oqrnxtoAabMgW3FbmYd3WBsYsAbV3iIKlDqYxcZlj2/20w4m2T
e+tWu7e9sNkTc/NndMUcTwhYXJRDOjsc6Clfwoylx3E5PDoCU6YaMKz09tD1oNUO9hLsImFd8Sd9
3yTutcfvPi0h9Gpp/7hoWCK+YC4hMbNfhmiJ9jiOeacrG16T+Ih3ezEnPEuU1NAVnCzXaPvEdY2O
65hNWX6RcMtLblN0sQaNeVUCn0uJusWTflXt1zJAISqw4tCA1BJ3FgmxvYOj7ytihG+FBZW5lOMy
H4GJB2NyWQPZcXqXH7Bw5GSKu19qQl6rjXaXXN8v2eZRmtdN1iZ3Yg4Q3Lhhvv5BT1D4EfG9vwyd
QWCqs64n+FyIWzAVNczx8aPSzN2RWPrAUeuV4pBOcXwzif+Resk/AV9xBZzplxBP7DqSFcCQDgYn
Rjhw0cx4Cm2xOPpmRbfsVNbkzuxM6dGrsa6z38E8wLoPapTsL4mkD2HcEwWkMy4RsWxn4wNaSVdW
QIpaO3tKGHNjEXfLNnG0ASz7ApelnueR8g0J/uEG2z/eejpCh45VWW9oqDqJwVAZb1MWmXJTdaF5
8bnY9hF2OLGjvQepP4sACm+oY+mof4kabBJjDiG4ZkFnVmpdeLXOBwwkhT/882wcQ+BGafpF7WGe
ntswjGXO/LDxjSmRMS1t2EhlAtLIwCGW6yTqIZTajUxjlTJfhNl6wxFOQWoun7AONqDgAgoZ8aIt
bGP5Lqfn1D/3i63ZOJa5/HXqJusfW7gd3ZzggXLPjsHSfRfh20bsR7RwAWgK0b7xJvmC0kmM3yDs
PinkkBlEAmIz3Z9W4EEFdFjwlBxoGegCqTO1tqOMpLwCXHNyK6jF0wPYhCEXOBIdaJhhx5TvUJD7
LINrfKnG/dt2VmUDPbA7937EqjcqJBdbltXLPeF56d5dt0td+shz5kXQ7uzSN9cRSCnzOUm41SaT
0g4fwaWPvq2Wmqs1GrDO/bJVomH5W9gjj2x+rqaERM7R63djbo+mdykxUtZab5rZWaro44ByeGSp
rliBuNnb06mA5HnRAI7mpjxZV2wAhVvWoxtLC2vXXOSvcuS0OxjIi5wVH8JnX5kt+bFoI31CRIhW
hBPOJSlBmOiR83kKFadQvLAswa3OPjYeLNg3yMpVz3p/McM5Rz+Yp7cdaHsE0Tp3eSCGIfYmpYZE
O5oaIbaoRVzy7cx8nPvpjW/mQ3kQWNJilq9FOM6NSQn9SIjxcxQRqqUKtrJJOBQLqn4mewu1QeT7
RBr9KaIeO5sTuhfYVLFEqpy9winO5lYwXVoJjBDD2ABt3cBhVBOjRZxbWtjfhfqqmyv/e7lrVTDG
Pk1AIiE5eY9yLM4x6faIMPnxMYOvuIIuhJiBDQj5FrMVwnX5wUuo/sEm7nTytbX+CPvOObAxcAIt
q+bP2qpz6vHkHkL37xEzoEE3qlfLdgj1XZV8/Pr+P78J397mlRZ3ElQF3wbSFZtussm3ruwk5zFh
qtGWqbRu/F05qFUW5wwdi5K1ELp6HMZo/MyT+uMqOHoLV1O649BXUhLvwNITXpg8RvWM7hV0Vtk5
elxqw6jHj1VtvwCUF3UDWwK7bPPCN6qTy0+Nt90VT/fvyoKBvVXkpwmla87J2NMiIKRUCrbqb25+
LiTOu0DWQ2J32SdroHae7C9bekg/LbGgTdowfp6UUFAdafyXMOKxmflnJdcMQOLZuZtbIM2uK9aY
Hzw+pv+VT50ECp6NyRQ4B8xfP3HkntHqFXZ7aOefVYGkQyMZC1O9ln/xZaOrLw2ZsqyoEPgILGBk
GA5EJkUOtq2DNNTfH63yYvULTSw1Hnuep9sk58M5+Qu6lVrjh2RIaMB53dsgznVzK3nIPfSfLSrl
jsEwAazMaqALBvLMa6Z7T6Cnc0FAbQZiNChYvPJnT3zHO4hIUeWBIY5gBLw+F7BC2EGETUrzt6Zh
SqU+WBa7iwmCN0nImpgy6ByQhj86XFLY7OK35Vp8033Az7X7BsDrvKwVzE7hQXn5OgE2K4sUff/B
6ttCRIhaPmE74mwnj3Niw2/Pp1qwkMNQeNL7Je7qzkvm8nf+WFnzGVAGnokzpBYpByI8gwfqPXIc
ME2N46g5EjGGW4e7fhZ20fP1GeVjRuA8+43WBcaR0MjFZGyL9iVAix+lAEOsLNWm4DwdqX/VA+bz
u1b2utFTQCtD8QY2uYHrct0ikBLmVd/98C9L7nhVXu2O6wR5zIY8YRxuw65QHJURXb8uzycOvEa1
Wk4dYnWigFod/db2C4+51LnlBW/qCTWDRMZ0e5asYLjrske5sg2SIffmAkpuZlNyJiw7dYSi1rve
jegQM8ea2zPZptyJjaoXAabE+2uRSjsAkcZu3kueVVq+VzYEI1DhepfDLgMTcrBwbdCgkEocC8wW
IQeQ/h5P6YVC5Si0UT7aRQH2tfxFs1wgZ3yUTip3w1ItewifdCqXP5WE/G4lrYhE6kWT1H+OiSf4
xix+3hYOOPLZLIQ7Vqmhbcw5ONHlrvCGd46R9eg/y94vvnFtQzS78BU8aTeRh29w2fouKGQ0rax9
bcZqMXp+NoHAF2T7prYVXaDYqsq8NbU8K+l6UIpTkyMbjnIdz2GXvEclzHpkJOFNcHzYmhXx+JwD
qZEpoG+vz32vl5JpGw/K4RrNMA/PDFbJsR3yINAV6jJpHzM9vVCMq4eDXDihpnnFUZuY4VLlxt0w
4NRR57gpiUwoNe9aB+AQ7IAvY0Z4G2qQjPTizaPAPVBJvr2+fJO0uGOmA/2E533XV8r23BMtTJjL
8HrfTgwb/rhJ2/HMGZWE/m/TlZ1R8MfNqvPoz6hwINzIoUL7uEzgfqrJ+X7JykpJ46F6JVZ6O08n
bOqjinNZc65kIAd7RtWyKpe4fdhJccdk+sXlpvDz485PJ+vCzdbF/DgnfhX7krZfrpFggA4PY1wC
mVaJ4m7ClDjSvbzUDEcMoK/40nTm5jVTu0TJj6k6TeksiHYXMC+lFJo3ErSIj4G+Jsalf7qbdhiu
8K0C/BbrOXuXL6qs4RmbZozZpZ2hBtPVwIx1LzXubQqJNTteJYjtHbNSBhKedUdEGXgVJYqQvVes
4pj+VJE9PQtmkhOSZKm0ciqPd1S/ZJdAMR3/pQ+wvEFmfsHDV4X49e3Ukr/P9hDhFRPk0Y556bQ6
lkcdY1AaaX7WP7rUVFDx/fdJa3v3NLzpODC53ues5X961oejQBJattVzND4SdKd3jHZ8hvJrGVSX
EmpCgKJPcs+mYJP66Ttt6J+Zza37z18YdzWrpyfx8PSBoU0F4e5Zy1vtOdcCsjxktS+R6h8ZwW7b
7Y9nOnbekAca/bQQ5BQzJPDfotMaFHX4Ju+toqLuq8hBdtQIftyDziSRrK7ei+MYaHPMfCW5DUH1
1LAZSBF2Oo+AXswi7PPwj/lBD3Om4h7Z8ITfEeSqyqBDu7peZzK+TD/32oPz5oVMfys0e5Z8sA0R
STjn97sF1Y9QTD1qN24xk0AOYxXce9uhrEO3hBMP78fjFnJcE7MgjNN2V+ITuuwL8lYbMMpyXyHF
qqwMxJwG1g8+GQsYGCjNpQGHNDIHV4j3PO6ukGaVR8TPeYmpOaQSfjmkMlvLXv0HyGW4D2i+eQPN
MGakIpHjL0VfyR/x86Jzr4JvIa/SznPJ5M2DEh0XllsVYQcUfcHZ+RfnwdhQEOXWdCYIoygJJWmR
W99DAeqhNhm+41JNvwB7WFyrVGOE9FrZdB1S5rNuEdyEQQnigRnEw8rim7DzwaPiDuzwPNI24EbL
hvOWl3TMPrbeSiZJwiH9op6eQM+NYFF3Y9jhpsOkwCXaIfC2aFkCKI1s8gICYgKUznCdElv8NcCL
9zl0t7ufLXvOcL+6fCHNMMJe1emo2WjxUbaM1HhPNg4ZDC3aA85gTRvVwg6BjdLSGIuCvW+/RPKD
6bS8D8f4tL1BGMR8w7th09XVS0v7kl6xcGIbj5a1hbcWoaOarUsSrv7e8n97NC/qD2s3iInA8+lo
KYbFD8DaGrs7bDl90W8tEfMk3IE3pY8nu0KcXsfDL0Y9zWmpsgWybXxuA7R/Bnt9dJ4qBcDVUHff
IxT5qapOnvne3zOt1cdP3IHhJGJOyo/S4uuRD8h+3z0kP4nSr/oPt98vMD0PIjKG6Btsfktj0xJm
JuWcHIJ9vx5Ty08DwasVKRziqcGx39PZ61dWi3msd14pnFcq9g2GkCxntkNvkXuV8ZaV4mgyceW1
/olV8qLMbUPLgA2sBE6HXsjG9x7IwUUNHEE6py/GClrFBtNPEIp3GwHElKujTWZEO24F56h2zzKq
Kb4lQ1vW3CEP6llvEEui8DKwBY2qRjFNBzUavPgHsWUQpFN/xP7emonGja9x1zZnbHNMzinBHWM4
1gEyx0CJYe3ZvAyqiyt5P4SUzOlTKpL/+V8RVAxrlxtQSBQUFWROpmmdDn5uItpuDlNhEIHXjbfP
Jh7LaPmHA4RJtqQy+jS6+TMQ+fPfqRD6t1yvVx8FIWAQ1QdkNP37xyR448/p6fVezaMHAFpcD0w8
XmNgXa1ToLvrswP2AEkvjNCIPNOslxaBZlcyNFKImyALdsYi4Y/xLrOk7ad8461CgJ1a6977h0Yn
jemF7JBpYq+zJPuqbZnK4Jwmjv0yDrLnzRz3NtYdwoDD4jRqnyjKdpfXYAz0OwCjntovHaLq1wHU
R5b0ctlHP6gJ3DiDbkDst14SOMe93x5sorvsK82PdtcmVxaZ1U2KW2mTFSr3zD8g0isVTNMeVIeO
VMkKgr9FtZBBIr3QQOmtnBf1FZH4UGQRyHL0LVDA9u30jnjLm4s6iHBoIT9fGcIEFu7NoECT2EZp
oBAsjlMwecq1RhiYtcjUdN5+xY2Jgw1yW/lkde9XdZCc41keIjcNYJFls+dS7Js9peoKtqq4SaOy
h9liMHnCD9AMOsDyjTJ1g7SuajqlrCM20TqFhUrSTLDsqZFgaDxrT/Tm/Ub/2hlAvPgx0t3k3s92
hneVj4t16YmSzBzNi6beW8sOqX0i1CYXGpMWGSkvFGGftIgN+10YhphTVPVQEKhdkF+z8S9URhQj
4aSjr/qWrvbx248+YxMs9Q3qob+LlxhYf7i0DMfuXJ8M05j28a0G//rAAX8+XwrQLAxbOz+Nv7uf
5XEpZ7vr0yW/86gyohF1/+Ww80FwgdLDcXFthn0fpweGRzPY3rmz12xCMJWlrixsXk5Ao8DxVsId
jMnUA5JbZl/2kXxAEI043S3p8ZCayYlda48WIwT6fKNsKMxizlt3fVLFD7RcCALUsAaaYVacnNLW
iLJiMjx44GYUG3wWBqY2PDFWIJo+YyD2il/e7HW8aga0XzLZyMG4q6RPEJjTExSJ9ykEtVhurP5c
8faFm4XgK7ckf++uv3GokwUd62Jd0kPd0pCDbRqy3OTnkJvQRUOUnamLf91abuQAvnhcWP6c7G5e
3Aagtq5EfeIl7J0RQC2SZJkJMb0uSO9wtLMLX4m66Zkzg9nhKNWoa35u/JxUfPpbCVrdT/KEmI2X
IOmyOISdyFOYVenhaxZSj4YjntOJCaPSNSsr7w4tmgt3PYROeGsuFVymHOlUPQmO/E2M0F4Np8Cc
tCPVVkM3ofbxtC39cRVsSb6TBJShVcst0okwRpgaci1mqj7GHMTog7PchWzFZBj/xjWt8evQ6/Df
9SisnIVF0cG129/WDSqddBMN1cCo7tDuQOQXS9bxrtBrgQfGYgWSIar4WbEnfNZCJpbXUlCdgBt+
1AjwAflbiYDvw3mVfKS8+39uENdI9yf7qe0ky2J9G4XiGI8FB8iNLYs0LLduS5I/+FMiHA/0otfg
lgN9U16Db+Z78F4hy92JLW3DZBH318sHL3n6958PyxNLT91T/RnNvgut06MQ9XK3Asmm7QbmBApG
fSYAB6ALCQkt4IpGrBt7ehNdC7OMyJB0oH7JsJ2JsBg8/DVgO+Mt2fpy0L0MDVb0AL2hLdwWNiLG
TwHUfR9ZpHFQei8BEQJbiZFsYFEsc8MTbXYAD0eRaJYUdO6TQP55N6AKtQxA3DAEXQxL8A==
`pragma protect end_protected
