// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cT4DuTaxQrLoQyK0Ltc/h4sTmZ/qanQRZ62VPKOHeDt4bk8FxCCEgyGx6qKVXhbd
zwom6S0wYYbRj/vQHb1ufOk2d7TPm4IptL84FUHTzCgmDZdQk6c6dZlfHNGh2eD5
93OaT/1Sp8lDxUrhUt8HTFKo/keEBKtyrhKvdbFpJVQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3120)
3MPTV8NfRuCSnUVD5eQ9xEPOOOJjKP6UVuhuSlW3LY/gIIiFHiMh0r+WnERSEviu
GcQYpvZiq8pYAqKVFkN5FTkrax1BVUXGx1hl7IiuzjvrmTwN61WqlDhIqOp6943H
4kUy8z7TKHftD4QaljfvjuyorAUfTmkswSojwuYdAwK6m4+alRY+m1+doS17nPaU
uQTAWeDsxQRpMCBP6Mx4S2Ltj3Vjbywm0J59WIekirPbCiF3eoUGjgCmd09VWfnt
96fvuo1jOYmkc9Ob9+WxjWwwpmebj7Vj/Tle8n6K2pTFg1DDwqAKUZ4ig1ZKbRIE
OW9cGU4ZEEyp7jU0p48mPXEHbZj+0d39jomUmkObUtx0wIAcUJpFLl23B4JD2qAC
V2x+MWZHFSaKLUA3W7G35uPfWhwG2s4H59ZasmqbAJT/Ext9pjaQZ9SY8ytN1MKN
PmxXO4Q+MFb8rfGjuySpP02XJsLRjC0AyS9uJO6zCuUVVSap43hsn0mHzLb9MHk9
7ZEMaAVmedn26EXP+OfDaVE3nRKx0DsGYPuYvLfr1hGfsM8lJXep7do9MWpbn/9r
7xUqBrQVqRkjdnpYjJn+mbV9To/snYzdOGd5dbpoGpYPGxYUmJWWGDq5rxd2zkZX
KV3QqfE/1xIDnD6o3xnLLkN4EA4txAGLeS/H4MdbQmD5h0BXCtP/7MCoNZXy2lCq
rZseLBhcNepnLqdor+0UFDAS+pOOaRJFfr0Ao0vm1Q/WFwIUX2v6fewMV1Re4LXu
lrJPGRd841eTcFJ1qq3CQ3MsnKVR5EPzRJDhXblb1SbrmIiZTqnCWF38Y1IhVG5L
NKahuaXZXOy409j9aEEfbJRQm0WdjbQUqCUyoafOzSfOwxAyqpQ4Ki/e+YHvg1IJ
HOwmsJF3pNAXLaUeuUGKwS48LBN2PNbS/W4PN+QgJu+nImDgYs3Ms5gWdEyXvU7I
+wUCwLyrBsLUZMdEK8cFYNhss9vk3z86vX2kJ6C8CV3GWeQIVZyJHqCdIW3VAhX5
dIRAAbv9AaE6FWFeHR8kEwcglRgd3u2EKXDtgt1KVFtk1gwc0lGJwSk2S9VrD1R9
70mjY0nLZhqKNwVtWCouThb/AsSjQlGXUFOI8Ywyvjlz6rCGsSOQLBeGaMTs7O1v
MGTtKIfRBtnyZMSl3Ts3IBXXKlzt7fbSZSpbeeRz3qb16Dvig00rgVyO9/dmf+HG
1C82/eDxK8tnfemMgTHqPNUCRnpvvyjxeSi/o0aOcRVauF2b4u/3rF1oTNHtLhB1
mUx8kyrcq5ik2efGu3212WN/XcW5s+WqDk8YqlGDaV8QJyQgue4VnEmg+mbFrDrW
K1gcb/oGsss+VAcJPyD4mc+E+gV4zrO+LOf5URAaIYtNMzUBK/LuGu7NlJ3222s/
uQA/cUe4pA4hdFzPUwv49oFBz3TjfRCSgA1tBnBwMJ0ElJ0uAdgo35GTsUxmwx2W
2SfSrqtjwgsQogoFmfNUq16/Kiq2dyBPNtuHwaMiUlokASyO8TP0fHDMZFftXduu
imo3pTyaikeVhm10Q9S7haUTXkxz6aIENvdQyQ9QBOwTQK1s/j904+ru0vaX6l3r
pTnqEuri4EeCmPkvYYcNjSfHIzQNRVApbTK/zWvAF7d+XmHXkBN60LfSHx84nc8H
ATiBZYhZd9o4U4bmv6hfiMXLQzN3/s9S0ljnGLdn5BqXTAummtGB8yd4KcGL7Xlm
rorSls//J4RIGlfkqOKx6W6oZafv6juP1DkAj40EQIQpqThQjcxjgejX2CqtmaLC
aHEfHS5x6EXoxOQbODsVbTwo3hTpgbE3ERZ8FKSA18kAQiWFoCaHJ1L8dHUVp06A
03hQ1PkyCSNLql6QelV12Ad3Ff16kPPMsqSDI+1CQwS17l75elxn2tgpF0J6AY8l
RrnEg47IXI4E75FvN/OrajuHVueiwg9kWYkO5p7RbfPFkXJCTRJPakOPqCSK29Br
OI7oIG3ga1SIDAmESqqEPGdP5ZBT3ZVEea3mQbOTLYquvBC8niZo1vS7G12Wuxd4
+rEc0fqABUUHfb8wLPOoQdU+y9yCKTo8KrWVBpiBCR3vAm9SPsmnb0ObgB88f5++
FCoyiQsJtDuTaiY4HzH/v4XVNolSmWmubeDUZS/GLxeMLhvUMWzesnZPV7Y6ZusA
Npw8Ft1IEU7CGXYKrNN0V4/kVBzP4PMrySVGSxk8ze9llLaZupOp9cQzusFMCjGd
eDuwWgYK+vfCmMsIZ+aKdkdbHlSbtWUQSUY4wyignG/gEWdWGBDu0cmuRbBi5l7Y
sQwD7sPvJSlPlPQV4MNofeMMtAdQp3cPgnSeCnYFf4EUfS1LSob+FiXvkp8mDF8r
jFHE6Ja3Wl6+fYsL7C5lFXlwSH193bLcK7YffBHaTsB8SRCNsc/7Y5M3qxgX3VUT
iWg9pMyciQNzYuHKqAvBD/l0w3ewD/esuSi9jhle60YU0W8DSZupCHbpaL8kkI6A
mFWRlX6CmTkoJa/h6egXDOUxqHDifnnp2tPTWrskzuV9X1DLkKuOROCuO0voN1rV
/g2/yuYoguptZM6MSskjjroqzWHQZ5Ib35FymU1isD3EIglfSrjp7lzgNzc/yyFk
GW67Tw5I1ZXfQ01BalufBdUNjRSXra+VDTYWsEsWvmPDlQzDylDZowU19eB41s7m
3II2Ow7Xt3uxSe+sQtEpc3tuKCgsC8ogAJl7lofnBOLs35NVLsOJQacEUPfD3C4R
ZOMqlwgS9oDxMFZxD+uMU7nBL03QJy3L+aH2aCE+UzlTGEUw3IyDfM31NjH+VQXo
zJxmx3PKjt6gDGUpIsFFBrU/TNjFwpr9vH0FgIiRIMrnVVnZifU0tYZu4adtRWcp
G0s6nzAuR83tuPQpatNa1kkvwn3+sR+UNCkmwev6klJ4kIqYdFk4ow+7RKyLN7Kn
LbByIbVkpaHlz+3dABtdfRTSdWrG8TV8JWFk866EW4103J2F13NW+9CHOHLGYImr
Tm3r5XVZe6JGUXF2/z+B8/zrZnZlEPuASpgeE2eQbqZxh2ja2cSH/3HgUIU6Lcpp
ROEAU1a4Z+QoDM+glZc1edOsiXu6omytOjvshhemCP0EOwI6DG1MbCKmdOSMeAIm
yPvtpv3XJRtdTYh//+U/lYBTf2XFO8mZPAUBt9M87Jg4eHZ/xT0Dni526jbLhz7R
qYICnUIS78HIIoqUOdfNDDhxu5WiTP5hJe7uSRLXwXbiQ7w8HkIJ6jaeQnaE0Pfr
wt0prclmMFqzxhfj3wS/qq/1bCKtuWxu4XgI7nDjpIFVkfWUdxp2AyjATiuMGbuK
E+OqZUK9klNxV/elFV3t5VhGOFyYj/6QZYPa6DAdu2bLHgmbBKz48mSQGVz/OsLt
gxaU9UXC/nH2ackbcZIllEB9HFQl/Dll73xlm4QrndL62Xyk1v2L1hdypSrMi7xx
O9VtoEXqYl0UYzRalHYUixL/iNeR3WH+oATWP2xjoOPhvcyhuJHkl6sB8p6NEvLY
H34FUzNcJJo0yWoiq7V8qC+o7B8sL7tLZN0d6CZQAcilLNgV1lPraLRqR18jsBrp
Zu0ApR9AMbzV0dAyzAeOPqnHG0d2ph6malM+GgTzRNj2fdnxnhfBqJ5rHTf9JgfN
yH1FwS+TIAqOO18cD2ObnG/eu4hd3P9CsD2QV/GLm/g/iZjsydGHYaZM9UHUoOjL
+jRDOIDJOSAu0jtPLMY0ka5IsyUC9Ujio8AtkN0ErqnSZ7CbJ9y7mdtCl2q9yP5H
Ld9Zox5u6rfoZmfUwW9yStYqyUkYAr91CSK1nFh5FMNzfB480t2uCaRQQ/ZnPf4Q
jEhpA8O21mr2xVlsrntPvdlEZbI4oIewVGw6Gfys3OEwvuwoaWcvN5DpB5C3zJ/G
guNf21QIqLPP0JzcIFFLAqFnbkFwJv+Xvdas+9LQTu9rnawqboQVp6UCo5Fbydnw
Kk34Az77K7LTaKmkApXSA2gX+cSyay/8YsSB+3Rb4y/iVvr22ez/DiePUSQjPq71
LWVe6NImbfYQztRyPihDlo4pKUAu8RsoOhmSNLVX9nENm+ZTgQ2pggecO+Co4bDs
B+J7Nep+lmvacbkXDJrcIkxC9NBmu4ktBx49s+Aqd5gvyoYUb3Aco49d7iuAqoB0
`pragma protect end_protected
