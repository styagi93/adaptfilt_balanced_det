-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bA892ZriLejgkhjey05ZYe6eIZRSXJhwtiDtU/4BiJGJumF71yaKb6S/sCsP5VH4e+vlqN4zOexg
6ijAdykW8fUBPHSFzDT8IC2v+0WKdjSJIWh+l8O7DSedCBNfd1+UdRtjbRsEur+gGx05a704x01y
ZumFS9EC3DC82T0O5pB/HIgcV9uJEUKWPJSVqDnyV3WMOOIJzgXW8kvZpbezRb2xjXn/Z3WhNBxq
8uAU2hsOKPTZhoM/bODE1u+O14oYf4AaPXDaOxtYnQS3Ied5sxUglQrH2zaAV1XyeXBzvCHl4sfJ
1Tr9fmAoNrdov50AAxvcpwHVhmnadFP3C8KIWA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7008)
`protect data_block
hUg64FerX5377BiQAYPdexZ5z2HSOaNvgGkWqhLw4aELX4y3/JhAAfCKSzkAQava3GEVQd8actWz
oKaQvwJLjlnCW6Ykc8EQq2HzmEA5sBLJXA/p60ouFzdK4VQ8jcUKWEqikBMGb1ke+h/C7Ejy0IeT
cw7E4dynNagjU55AdE2QtBVGXp0ik4mjKYt8KSwM6ugKxscni6qA/two7bywaX3CJU5qPB1ElQ2v
4ZdpKfZlA2tAA8BBHA5fotk19CVvv88sSMf4vb+y2Srud/m11W7UEs88EQhOo/JT3Tmr5cFEhVEm
rXvo7N/BmsfA9/yO0Gv3PLT0QWBvoP5BKCoCNI23BgRuoCDq4u3Sfxxo7VMOvoE4zkLREKhD1pmE
A0wruqCxMYhsULPhjEJjKvwL2zCNansrfq7TMJOjgyhkvaqRMujsBwFES6JY0XoLjjuhqlzIJodT
8Z481LzBoyefnJmm8gMwfbkF/kGC62dlte0ZIvqOl514JuSinPbQFdzsAmtQ0fwwClorUM26fwDl
qL147TW03iTwC7A+1qdqDcFyibZqG0P5RhZb6afAIQ+sKq0TL+hsjyvaU1cinY48xfCKsgG18WVv
x6T6U4T0StuiVG3+AguMVoH+Frr/a+qnRyK4OqUlAEBVw4dmh48dnBJUcSprXPPXvCguf2HFQpil
m1Xtm4iuH6eS77Ox/CTj+ZtMMXmMzjEP1duumvfIevKHjNLwvYSYP6K+JWpj5IfVCpss00RkpwVw
QOyYnyX2TrPxHzftDKbZ60flukVBhRJykP0YOsbkQRYrmO+i4HjODuCIwEAuMtr4MJU+EjfB/qkU
94vY5ovAL10Zrd72IGt2qU3DLeM44lwxH0kEyz1OuaX5KJwhKJjzWodVf9hGpt3BlQKfUYGFMIYn
MunNNcAPtc77iNtoHcKybudVj3FmWFZwfwOF0/N2+KAbVUlYqc/0jcC8NrxCsyTS78DvGrCgZ+Db
7cHOq4uPP+X4VelG5NWMIzkdgvhYJJ1xMdhn0NnzNs2z3yVaab0kaJ82hoM1/PQb16drbvnG1V/5
uLK5twHWQFA+UcP5wbD+fea3ZAjN8hJNJIrLQSsspM0TSOHy0+xa3TtzYQfAwtno05iqQZ3E0nqa
I3nrRIutgH00rTfKAOWkMyFTD4OTiW3ZuAJ9hwMxnrlrpEg56blRo4sV4Z+Ku6JZyoEwp1t+iSc2
DkdusR4qG3Cicobf/QIyq8CGVgdc+eLgV2o2t+nFAlCvh+o9JfxFOkc1XK20QPZfaScE8DEKAkLT
GwzYF4SjRKztyy1rowv/NH0Ku8AvJqMuQasb/O7vz6ow76q8z9fvptRnzyA9OETqfqNmwjyjF6NX
OFE3daKkNXrMXqSRcSs7j/42JWwD2m78WlzmAbUrpOmZvtQIsrTsLXE6VJ5nYZpCyPtKKlMvLg7F
1ijiTXk5Lnbn/T4j1DjUPM3+po1saq2LE6iPcBGeIG7SaWBud8OGU2chbTsn9JFY3VqP44WB6ay3
GK+1eHS9vLzGcFJcYlJ/yprfOp2B7aH9o/fuo2eXmaaZRohC+FtLWme6kdtnKKutRC+RiadXR9v4
MfLoimmqgdm/jUZ448cax/m4sj6AjPqI0t4sy6xRIxSOwPNFAhn4VpqfrQ1TdcHAcfV1HYVYnMIV
fh28Zk6oZNUY6s06kcmsIOuyIEuH56BkY4StneoCWvJgzRpCNOeHqHJfyfpJauecqi2nKu3pk+be
e0EvKbDojEEnyNOwX6OtI7/h2/6iycdqF57sNMk+uTotD5vCeNAQo8YZORYclf07g9OhGxQWFAN5
/P0mzKcryjvULUgDJ00NE+549gFyvc34VUVce93NDAu2RSlPJXf4/zJ2eTSJrKhSQtwCasZoF+Nz
s+cGLNbPmArhPRY4V24U31SuTTM0GoTEXodcxnIlyxdporKf5FIrRWme5ReKxOlNHN+bzRX6HEQU
wdczAlzXZ3OJCnX/mIhA4e8OtvvcFKB16NG1B1sEutlwT8GWmOIyWw3M8OVKH7qWZ3DPO5Jvgxd+
wdd2ZHNlnPoOZpCT/FfJh0xzrPxv0VYSSNRfI773xOFvoeQfQ0MPFxRUCfbjbZbtT8n+8dEhaxx1
f4QZLXkSjQeYLpBJn/ksbtQjW3ZTFHHryYTGn6wPdAAp2mpUgdRRZLDxMI9viCPGHqkRFoNBeKT4
Ivo/1lPVgG8ObVRj/TK1WmUCyoUMzJxu4bz+FjnRt7Ykni81upr7imAF5KXOzA+egp2a4B4PJGDB
V5Gu3Ew2wjkxgVNcawIj8P3BgyXI60Dx69CKtW+e5X52EOiYshduIx7TQKpsOe9A2kce9ozTZouC
1/pqozZ61HpCPhoMb80sFw9H2vPBjNU2d3VVifNQoAUalF2L7XHyxgVERUn9q+dBzU4eDlepxVKx
On3ahNIK+tXwfFR/zx+rVE4cRyfH/sxLtAKAg75heCVORsy3SUpqS34eDl6fneFhFInotLDtiD6u
QYoBUoNB2PJe5jtWAYKeWi9M3XDFPsE4h2lYfKdjV43bvICJx8xS5mW3p5hMift25RpDGxusXp1a
rPX36gTLPTvUasukP301NPKC56mrsHaLrjvD8fToWTKZ2I2LdfOolLLBtKio2GMTHrSq6wrNbrQD
ja/veRLgRdQm8CODfJnoMXooj+vTdh+5oMSD6/MwimQInOT45pd/e/2tek79IFG2gb+H8HY+rsKg
78+yZwxk0eyLD2KytWVJRsf4jQEWUBFdajrT0+cL2lLwlHxMKNUH0vKFextX3a9qjGujnWpLfCPm
ioRisAecEm7khZFzk1KlSTYWowQTFhKqgF6XEnkqpa05rWZURl37Lj0gSrUj1lyCHjZJgNECEiP/
m4t0QI9MD1ueikkujNGrLYGNAe8r1XlIgXZV7wnI7DSoPpI9f6U+U1W4wFR9NMVGu/cu+VTqfuCO
FomtkK2R8U2W0MP/JQxQeQrXtjKRhOMUP/hoqkpjo3xsMBOMLeZvl1EQbdYlP1OCDxD4vESiu1lK
2Bt0C3rET/+kK9vmJg9wzC1VozKOovPCRg4mQ3kaWgF8ZlvMQU+NNQZrzrTBlPzutk8Hzd+MeIiY
6nxtFmXeSlAZY8wYaY9qqcHhrop4IwpojJqqgwrq91UD+Igj4lvb+edVaoglLOChjWZIhZyUou9h
HJyNfQg5dU/QUwnwYIRbKeS6AixcEeDNQW1boMpzAuTKjh+CMucmKshSOVzLzXG/hsfY2xFVlI9v
njGz0nvN8x9oIhFngAjh3OTANA+7KwQ0HAGmcdrdHNoxk/o7VZgep31F1x5TWMK/LH2YbyNAsdIO
RTIGpVyWRoJm7vhH6zyAucqkdIOA6pcEle4qS9qpRaEAftxzjEMjMe0G8+D4iBaf2kloNqbQEu3x
msdaadWND1Hr12izwL29iwrMn/kd/hfqdSPfVrs7l2jXXhgcAXGfw2+/eF8lVzhLxzERd3dfce/m
MnyZUe6KHkNCPj0ZqVF3lRBZqECge1tFl4YgvB0tGKhBLQIyH7AErIwecEvBeFL1RSSbZUJAZZqu
WVYjAS135xec1Fh7gcXCOyN5FP6yQRxADKhR4hlfHbmx/Qt3+WxNNOhkHpjvmX16RR8W4oEmkR4a
4kJRpIpOnK3/WE+/2hOvCtgrPDK1hK336C0/I+mPw1n+HVqRJogdBdxT9WhBh4pXRa0FnA14fxAe
YaN9ijSNbjc///ZknxNMt4LFPoDwQkOZk+LtJUJoaVkAxmu7UtOJwYSno2zcJUTXBudS04Ko6EEz
yrv/rTxxKYBnwhGahXOx1R4wY3hcXG1w7+9hLdW9Uoh9N0Z6YihDBPvFqp4QJX7wy3VTsyEB965S
XiLyaBe4PsAE1d4fzhBerfguZQvgU1oRh/SueJfq5O2hrULRk+MjEkBO1Cv8SyB8VFrkKEEQT+ga
kza22tahkEuUXZmIrNEZ6drFjFQR6E7TKbB2N8jPvWqRIkI7jg0awR1C53gpnfZlQgNT+TDhSHa4
jXXk75sr3Pdx2P+K0UVtJN99fb5wIve7WeBR8vrAfPgsv1upoq/YOOrGf6F6EJ7di1k5HZRyyTyV
L87e/5SuigFkgiVh5fdEEJg05TLpN9bMLzfIt6krhGN4vVfKMDBUi4diNiKOW/fhH42eZyYub8ut
N6KAwCd+Tcg1z7WDpOruZIu6LO+HzcDfWCQEzJbMmwQCDcs/VpLJgTb8pZeYgBSWM90PrQJYI0Yj
ZaF2YSyEqEZwhoZVRj8vUZ7M3XuR0XebrOWAydEhIxHqF1moNxHcIxzZOHtgRJZOm/YDd/4vO9Xj
t16Hw25AL1XqcrahGT4ZHs87AmyLK/kpJ1P5qCIf9cNpbivRKGDbs0Rm/JEak0O4ZJNYXok8Vd1L
LjHQ1V8W3lQqBchISnTW+jZT2k9i3/k73ZEaLyDWaRQ2l3QXV2WoqdTRtSO7TpwnNRD/pL3VS9vq
yzLmmGbbS6gWOAU8uKv+28fK5sURBxyXfDgTyb3YJCWlMkM6gcRcCoOchUeuOlmMqxCgqmBLMRp3
oWz5Tg4wpAqBDKlQ8orGH2EdYc6Bm/fnzg5IdmWrZP4Mer4GZIRi99FFlHelQbZHXYLJhfNxm3V3
57hzWsKNxzng71vdYe0U/ILhIhRUqllqA+H7rcB2ncOgQ0nnKjxl6NbU083kEB/7a/J5VfZt1ZVa
JhjDWUIcpJstNoSBbD7JarLy6cLAHehxILFtRAEQslN9ENuLugihnFL+vBFRdi+vrNhUbQxLVRo6
H0Cu8I8rxVAgvcBT8jxFPBjYZMNpkGJL6EtJQZvPkE470P2n44e/o+owQhx+0X15mffVxQ962RzK
5FIzEEGe0FE4AHbusNJN91ZIiBf5a2c7YGy6yGkeFlMFDDMVedDLOPUJWvsB9W3CpwQPN8tIFFLh
iURa1BRlQlcS+Ynw5X1kvGr2OTpUB6OuuhFRT1bdqJaRv7JQ+PAxZ8vbTVxpywLR9+sZ0WUpGTU4
eJA+dtxMGeM0q6aNI6tOYblEglMzYkEylArYTP9of7lUT6RobGUQum8Kh3dF8t++5b3mOVym1D0T
EGsObDtCwXX7FVJnQnpl+1raUp7UL6TJA3BhrToRiKqQhIhdQQeeaNrsROqgcOut531GYoQWYlxN
4N1rYcoCs2hsS1Q9u9J3Gp/r5idkCI7dbysv+M5pQtfOX3xdS0LXeU84Oc9YtVCORhdjHQfP8HjR
bWBw4WimOEpwtx7miQyvZii+fJlfHjtH0jQW0JK95WUgf+Xlk/1JAhzDYs2r5i5H5uAXD61pIVda
cqrfnCfULrZGPtXb3H1Z4vajWLaj9BW29R4ENxVEszt+qu1WDg3nHMTj9w0PTV3AyBjK85+6kyv9
CsghKQJaHg3Ws67P9EFIYwUkK94EwAKo/SlmsxD4q4aiQ56zx1yEoBcAcZSl0KKm03S/D4gdUNia
QSzztC+xzj7LnxLuZPr5+KKzEzGX/wnp4AvIYSR4A5cw5q1pdhzfnWX/JR9b6uw8QcaCYR0u9E2E
PseFuocR+6udjZefqJ4gBsD4xL5kv/POAeGmN9zvjBK65G+e84vMRNFXW/NOt3MSMctjPe+Lk9tB
Hk3vlq0TrdO3I4/b0bCjrVLmo/3bXBaLbkWO6rBKZBi0yZdZHNIFaU4dygCqYhLKmRvWeZ1+mWmy
qTI6TXGlnau+SkXVcroI7Zz3DtS2eKQMcOuvWh4wy8SVZ0IXe/Re3Pjaz8s+FFJEx91Z0x0qC7Fk
+Srcn0Al37C0Gg8j2MDaXl8NzcLjpHb00cPXzT1QbVQzgOV5QARVf7HGosvsVZtzJXePDjurdnzV
Ch3ZuD0mF9YSql9hmeHlVcO3mGdMNvYAqhPy1Xa/7BtgoQuOPvE526w3dPnHQQZlpe4vDhXDoypJ
r3wWk13b6ba9ldjW8i1aw766ORCO462hqioB2US/He/XNAKi5LM0tg0OGt8q/PgUIyyF6yS4haJM
HYSA1bBby081CLKkiwpWu/6TL7cYpZpF5XHeIWcVHAsgd1sz1qYWzCMOXkYJUnOB15JcQ/f6zZJ4
K+8Y82F2F6C49mG5Uc2cjoQvUbZadqne62+TnLdEDkAdfSQQdC7M00LB8I73DvPKnd4fs0qBwhAX
QaXKtjvNGSnzfF+GTzSpgNn+GOVsBBiEfgfaV+u141JElmzEJ8DqF+5rzhf1D8ww6K3sdTB+iFDV
/W744Ehmk3fTrwmw9Hi/QRQl6R13kUXKRmSfzirgI4Jtsq0ByPKCxaokKAqOqBOtob928P29Xm/t
mO6zxrTMDevEy1NdQkvQy7zMWF9oL4Lo78f/i3ku7G/P47sChlYx29lFP8jSVdkgQzqTF1qrJRIv
UNx9mjjO+Sigz/2HCqq6h1RgY3XakTxMK9MMMinPAk2DbiDaMlRexYfp1bb83X78NpZw6J/Wafdj
nFregSm4AUpA91QzvT/o2UQ7UPAB9ZEhWodjneVdBokXhaFn6LYeZeNzWU/T+IszahZtwxv+moBV
mbSxGDvT50gQm3M0pUb5dPTjYNeeHy6OWuvqVHqpgBXT7XVWzDfixHd1P5CYmSiDkvM88kkNlouL
6wEC4ZWw8xho5zYM+2CGwrq1GOrUGXdApoBjGIeqV8ZFCh4CFyVNctmzMoj6HtoCa0q3PNaVptkA
eDgOeJA/c5/xYBG/iw6qOcGUGpTY3Z81QzgaYJC9QMzaTUS8MTOa/N0b6ZOC4Wmb2MQf/yvAmRun
JuxDF+M2yNrzR9YQTQZLK83TQzEvN6xbsK7bv4mpqPIFwpp/taAzJR3nhIlTDTD8US8UF+dCb4LR
X1N4RT7r0i6MVkeGoB82CdPK44CDQ2nDjyRRJJ6nXeYMckgTaSNMyKG6z3etVNwJk8CxobhmJDNT
7bBDn+3yzS8+/j7eKix4kCEj1w2XaR5C3yHpmv+sqPhC6FFRR3tZ9PJAX/CoXKRODmB4Jfx0DpB5
lxEd3cpyT7tT2qqsGHD5ADR6eeBY8mYG2uzAs9oV/dLg4aVhd8Y2Ij1p8SyIitOMJ1hei3kBXkgV
2oble2O+/jnVRTDxvI1rzherRNth7P8ZhD/M23tahQkq2UloAzkZB0cG1SIEc/p2cah0EsQV/6HP
VTRvsjS8jITuc1mnsbFdv1kdEz7FDgacs/UkPEKvwuCf623olAhqaKEDosJ5dNpG1iHMBNOCjCrs
rmxngt3bRW5oTlMYy7kjnmyJYImbMoToGP2jCkN8KWUSnUCfxp1YPK7bA/c/Xeq2z1uvSkn9sPGk
e6X4uBsgNMGAZJMycP8wg6svakJO6mc5SWoONbmvn//VE8P7QQwAcuzZxbC3E75HMmWybxca+VIl
74ZHQSPtK1qXZgwOPMlkAqU7k//TOCbBcT9SC3O4ZxD4p3kH+Q1mU3oseHsXjTlvbzEveMPx56EK
GC9ChATlr5ilwrW84/QaMGwGvSnYGPgOujIuciCE993R0bZUz7CGY0JRd1e6MAPOqLHiSnLKO5Ja
AOcgFoTz0LHOkneFCT9uk6dN+RHSuN9FdgotMVsZAW4K/22mMcRHjyFGKGozfNpmwsTbjdik8qz6
D/eKZc9UJ6xIc1Z/9TIFcH/yJOkzq6g6m3Zhom8zW+HexXz6ZzSbFJJlhla1UOb/Za09NDBUf6Cj
IPA+adWeOsGH5KCFyhyX9wnWF+qA07Zv8U9fXPt1EDkoY3PGM7TABkhVnuPbo/+mwx4iFzjaG6fF
i9pbwkpgzlHzPGfWNHyciAdju1PwgXumqszL4C0wQKzy4tgn7tyjA2FLJB5qnvT7DJfJYUqKeOs+
RjfFz6nCLhJ8R5BHzV6CIqshBefdZhqqTPxXwv3lFp4j+6QsWYBdVqRtuYgOSHwGa9WmNKaC3RbO
/BCeAf/dtJayrA7SU0Iv+g8bkwquFuH67ynTAj0hN2+mV8nm0/fI2A9eG7+NpxkgarIasnkzE14c
PbDF+Q1vjnyO5m4+Savu6ahw4LnfsxS0KbFl/dqpQAonvFeZ1mx6YdA7U9QgkoTrMqx0BXT7ohVl
s44XCYjo6dap3vclfdw0tArC9g98dh9sbo/BSpo1HEj4cuf2txz3sLB5wD2xHNI5n/bFDsrp4tYU
h0sH9TYT6BGbG93lezJ+KUojnpCit9biT03mxb81yYi/niWR0Mzef5yBJ0EtlCdpfzcnvJF9KogV
62BE1z4FyNckba6mgbdthr160Gm1h2DUAN3i95JGX9/4c1zo7Kb3x/ipH6PNS/UPrR/ndGmcGlib
fO4yXxg3nYmcIbp6c1J5+O64TcH65UJQZuvLkOLHBqavg17WC5W82c6eHaI7UX68TZhlZ9MZ5wDy
bVkQ+p20jl+ijNgP20+jw6AZ/Kxq82ImbWine9x50wqpzWPG+DP7+bg6+kVNlHpv/D290nQh/cZN
QQl4L8HQ33aJ7JdTN7ZC59mDfWJ8TF9k6KoIK7B8K9hi+35geFozHve43mMRFUpJLnbY4Q8f/35H
r8aXSwSJoLy622nZwJFaSHgdahuv7Du72D5FIY0eu+ZcuN+Me9A0ddh+FgqIuf79nWfwQ9Qz1MYI
FMo7ssLZ2F0TgPoR7uZjl4Nwh1jetPcOHr0Q/eOudnOfmdA+Q0uXvGK2dm4Pxgd+djsPoA4a+JI/
XEubMrje4wmQqAYtjxatYuN5uMGbUzBCWkRKUGhGXxPUcj21NsidIiFW+ePnL0flWciASG1a92Yx
CSg6+l9Fo7ebGDyCjV0AoEsUIGxalXtZ8HHUwmlYH9aFaSLdk7Qb1AZ4GFdjgDLgqEj04roFT7pU
vg+1OJ3UhheYMm8wv/cXroBp4IfaB33I7daDh+s3RX8/+rbml0lX9aBljYglkVhmD1AMEull8rsd
VDr78Ar+o0kdmZgO1XknsMObUdzKsI0H+UGEpHucg8PbE92uKxP6+0D/SL4mX8R5RKBu/DJj/hWv
if1SE8/N0o0Y8R9QsQPw3WpCsQ0bNOPVZPmKkwOyvFsYT3beV/MLokIdQXzXilkzfsnfSSuB/7wt
//TZMLdnrAiW3tCiiVsm5qKppNCOZGPSfpk0yxIGvv4HT15W4wgNZ604pfq5FRIjWFeMcFZ982sV
MyZgiv2e5ztWCdqAiYCQ+rC0rh5dhF7u9toJxW4cSncmZG8YUMm/mqLJ9cZn5k/StokTZJ+T+/OZ
40CxwDkERz6K0gTesjIPUfuW23GMDRwtFop56BT7UTB7GTprtyFB+m3fEmbbY7pZyhdM6YDbWpGx
5e/ljobxuclEDGBW1QIukfYKkoET9/pF0Ceu25jhbFTHjyuvnjjVGEqeYw+WcIG50V8xtHtL
`protect end_protected
