��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|ֱ�}�7r�v����ɤ�⑳���E䲭�	���/����E�9��eg|������v�(��	�%m��Ab�+'?�.�7y�y�U%(�g����Wn�-����[�:�i`�h*��,c����2� /6��Y�F}L��Cg�t���v�*��T�Ǹ���r`�@ת֢0�x�qy�6�~���؟d](�&Qʆ@��R�9G*���oXN˩x��������*b4��]M������נ�V6�HRɃ� 0� �[�l�.�w��}m�K](�@���9;���K��i��/_�l[�>�~hSæ�~k�d��x}����!����]�V��e�!�N�%,��/ր���3'(��P���Ⱥ��3�����Q;���f�\/[)z%N(1z=
����a��_��0����Y���Ԕ�"��X�������"_�u��s��ʭ^#,���6�vA��r�΢� �xY�����k����4z����<%(a�^G5M�Ł�z����L�>�k����@��l� iF��8��6��Lo-�94{&��f>˂���f�w_��[���3P酹�Ж��l8FudQ��|�e���'����r��࢛,�Ï�z 4�e&_W�>�@M�X�j]�G*x�!�mA�v�z�����.#��J��_��q�%y�&ƫ�p��w��<�}0�ۚ,��P��+�ڽ��I�	�l�ɈY��K'�/�d���_Gr�:������bm1��]�{!)Q`��y�y^ehj�s;޷��q��h��2�tS@P�Ez�^Zjn3�����w�#�Y�����w¥t*���*�{�]1�Oy��sD��y&�}�څ���1��q�����7�b>4�Z%���Xz�N�-nN�^2��Qw��|Ήӓ��*����:E��w��2��Y^ݪ�%���u�2�aW�b�.��L�܄��j�H۪��[��1iU��/�k��^��K�0-�Id�)��Ei�t<�B��X�bL"��Z���$B��"ύѯ��m͓�a�R�а/����6���U�sQ>�3��gVZŝv�M��j>�Y�7N�`j�8�G{(�1�:Ժ+��Z˦�VS�N4`��#�ެH&��NP4�g�U=����Viw.i�q�����Uie��ߍ���9kX,���-�;����:,.����2�����u�B�5��Q�̑�K��u�8���y@y+%���ӹa�*� =�e-��D/���yՓ�A�i�O�=nǵA1)%��VN"0�LQ@>�b�K7��(Re�;�f�Qvg�D]�ǅ�j�&U���%�D����o�D����j���T,v�g�]+ȟ��D\}�
���>O8��~�'o�i1o����Rs��W7�@dx��j�/-��`�_���d���@H��4�ͭ4�m�?r\�����$��z��7�Ҽ�0x;��e�4
�k���N�mMp��IO�P_л��_X�,"��NgL�[�s9��ϕ�����/Z��P7|��J�x6�I�F��d.��C!��|�}�/�S�.*C(<��X[%_�S�:
`usU��}��C�e�)/V@x_]�HGM
jR��W�]�p�@��XO��ܳ�zB���^=P85X�B�+�O�J�Zd�I��k�L�o6� �e.���G*�ҫ��_��8�+[��4�|$�[r�EHW�(#s��mz.ʐ����q H�F�� ��^��W����l��I�[E��� �7R+g�A�Wcj�p|x��6#p\ڡ<+��t{;�%��km��4����,�?֜�H(׉wm��r�H�z���ٙ���p=M>ɒ	�nK͈ 6<�^?E�G
Fה�,+ͧ��xl;}�Yv�Z9ٕ�>�u�GL�K'xN��x����ܟC*1����E��Wؽ��ϣ�h�O8��y�#�_�J��.c	���c[P�0 eC�y��4� �4d��%G����CaJ��]GVu�>g,D^����Kɮ�j�2W>�V�Iz}��8+.��Q^�0hB���$%� �>g�њ-CSu��6ϊW����&ںr��t	�0�J|����ؤ�O��q�6V�c��9R�+�C��m�������mGkyx��q�Z�\Q�{��>��C���9xc0҈A�jQj.�h��.{���8�=�,7���(�L^U�n��6),�آ��p�	>�i��!�}Z1� ��.7;�ŵ8��q��B��^a�5,B��E�9A�E�� HT�n��)AN�KA̍�f]���������r�K(��:��r�Z�	��S�.�VQ7u�,䲶�W}�\�H����u2R�y��;+A��ӽ��媭�!�u���p��R��Gc���Eb9�~:��h3��N�j�o��?��;��e�U��]��2���D_��k'7t_{nFڻ����A'�t݂/��C�R��G�Z�>���3Sz4��c�SO]A0|�ʺ��~�j�ji�C�L��=����G�N2�N}���(y+U���T�b�l�*�?D�7K������.��?�������zb��#kzWI����C��Ar b�'�S���u��i��JP�wgQ�T�K��5��Om�K�7�Y�����(|d�N՜{��V��x��m�_�o:Yb4�gq#�/��#�J_̂l̆��YF֧�q��K@��s�+K������\��UX0���߸�/�2��M��}�?Ƽ�ۨMƔW�Umy^S�J �����S����\,��FK��+P�XF��K%u�@)�T�WCb7����h�JB�\�>��0Ȼb+���;��]��F����]z��~���D��X_��ۀq�Kh����������h�JF*��"�ٺ��;�
ͩ��*\A����)s�;��.�������{f�oIh
n���OC�b�攋%���燨���Jǽ��|�q�cinV�8ĺ<�;(|�2%~�/��"i�YH�p.=�^���ĜE���蘉;M��}M?O���VB*�S}� �aI��:�J�!8Ƈ��[�}:�E�H\x*��,ȘM�����t"�^6}8��&���� ��L�+7��/�e�Q�/�NX�mm.�]�6b�g��J��l�,�g���U?
ր��0�9"{��C͢�U��U116��M����6N�P�,Dgp��.Ul��,]]����yhMRnÝq6�s�*-��X��!#b&�K/U`��7�ǔa�~�$��s�A�P��T
�|u�T/(��Zu�){��,������@"�+�u�L���t�B ������u��Pf�ƸE�;�쿯.�	�7���S�Bĭ�T���=�1�4�%�A�a����|�4|�/r�����P�VK�k�,���GܒǫNև0ZM���)Z�c�� b�08���vC��IIb�B��r����	�X&�?�q(~�ڗ���y��R��VR8�Y�0��kBF�ۙǏ�b�
���K�'���_1O9�`���m$Sr�\�j�0�1 r2�F�z[��6x<v�E�ċ��2�T�!��N~��t��.���R�eJŊӚ\��b	�w���.��p�-t=��гݔW���@�ˏ�<�R%P�Dgg�	�1��U]��0:�lv _�l����(0�O�w�Q�)��#y�О�v��#GOc֜���\Fk��G]�����g���z�쏟B׆{�����<W�xh���N����N�!2ǭ�,ڽ�%�A<�QO�8�+\��,a
�n�]�e9谠��]�����z���f�jۺ�����}VRchq/���[_z��Mm!n O*2�u�Q_�����+�x��6��4���U?�k4�7�Ƌ�^��d-�^x� Zf�9�Ң�'�0���`��AO�}�;e�L���6���W�v%��`��w3���x 3 �)�3�C�y�Qa������^F͵l��5S`�N/�����]�/v�R$"�����/m�bJ��Oc���.�,n?��%�^�m�{^�w�G�������S�A��PIM��!Z�	"{|�b�&Y!�9�m5\�t�D ���$��rc�����ԕ}hմ���
|�l��v٠�U�����	J���	�~�R�Y���u��8����Kurcmg
v��AN�^�B��R�������An��Ɂ�x#��b8����j�mK(nJ=B:�dI��=�!(L��8V$�����[��u������m� �1h�&e�' 7սx*����q=F����Z�c���-EhP�*�
s��"��Z�O�����X�
1QYPP�`��*N��l�pHm���S�߻�-��*����Z�aMr�/���.����Q��ChM��%]l�+�P7X(f�A��@�K�� ��e;!%S�H��	�Z�NB�i�A)^�
�Ng�!i�#�^V�7��2,�?J�G-����CX8�����j^u��hA�,�����'����$�ǜ�_Tz�Y$>	��y�/������������J8�S�mE� �E��3�j���X�x����$��X>��k������$���<K��Q���iM�,��f�k]N�s��>ꇾA �3�h��
,&�`���z�`:����I�lJ6�[Σ�qx�r�
.�a���t�n��Y���+��#iN5���e�|{���[��e�!G��IO!�>��:���S%`y����7�<ǚ}QZ���Ɯ��k�L��@`��OQ�!��S�ʧy�6KU|���Vzc���ծ:�h�yb�O)��U�������"�A��Μ8`.������A�g���.�:d��?~�W�H���<=��)�M��Z�&U(��E���#Z��ї�EW���ȗj�7k�R����%:,�0�f%�	b��{���<��^ĸBf�7~�ܭ��ZLV����S4��S�&h�VE��u�����g��V�ts>_XF�(��ZA�܂M�<0F��L��b��ם�wh\6_���^x�ⲳ(��vD~wܽ~�^�z;'�}럫�1m����Z����{m��I]���YLGIݯ�tN<�/��B#�	���a�ކ�Q�!u1��=��Y����xyuV�s�qj�/��ӯ�,C%�Zl3�+�E����s���niTA+kCKҲZx[�䝏^p�n.���4n1�DIH��pz0�/��q��R|�LK!
C�-�5���P�.�v��IB�#^�q���\�����M��k�b����O�\�m��B��l�嘚�tEJQ���Jg��:��v�2�&8j��%h
�
B?n )2�R��`Ń(�Q(��7<��ըJE?u���`��	��r�i��ړY�g��SR���W�ͥVg���������'��m��|�#��#��x�	_N޸�!�m\��U�\� m�r�,��@�t�챩i���m]>]�C��(�<�Ef�a;@kօ�!�K ��a��	�L��������O�?�Q$�1�>dT�.E�W��[ �`E���;,�9&G��޺oy-:��xO
?�y�� ���|�3��Y^���WU2��V������Lk�'#M�HВ/wkZ�e�}��K���'3�g��e��
��d�vR�UN�8���`T�m��]P����%&��7������R�ͦ����?��0Xs�r"���I�PQak�bT]{P�'2/7ȚБf�*�Fj"�@������%�>�4w�ݗͩF{�=]#�RJW�E�P~]�~<��c�v�?��.�I1IF����\�I�R��� �C7�L�s^x�&N۔R���UG@a�&�6�Qe���b0"㑹��(���,�,���oz
�z5�S�աz�T&���O���9/H ���96	1V oћ6@��V;�;���$>�����96tI
B�Ei��ʊ���O)�(F��o�+�&���iU�ֳTg|�+��/h�q��2bc��J�^�����\G�$�bܴ�W:X7-_��Z��>ѹ���?R��"�bl��w.`bq;���	�S&��V�y���ٞ,�D����*X)pmì"2���a���}$�`��c��L:���ߟ�H5q5R9���S���9ambk?\j���W��詂�n�(Df��j�n�`�ށ�Г�e��T3%b���Hl�-�g�Wz7��H��6Yl�kVB���B�@3������E=���9�1�Ø��C���ua��m'^��!^k��3������w4��l��F�u進�>��sV����dN��;>�-�s�-9�.�ⵘK��(~|��7:���<��Hq��߃��T��Ov"~f����S�G��"KBi�Ԍ��"��I�̾���