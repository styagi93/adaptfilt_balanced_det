��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,G�ss>ʂ���ܝ�%��mz����elD�h~�� �vx��Ӿ�����	��n�&���Y���f��o��s]]��ޠL��|SзZy$}d�	 ��Z!�dЎ�?�۹��F�_��ܱ�v׈�b�6��"��*ۊ�\�����J�UR�Z1W�{���ߡ��Y+|���P���4��
Z �2;$�/�&�K��E~-3�BB$�q�T�M��!&.�o��S�6޳�X�w
���dlt8��0��0Rc	7�3�
_/���Q�@-Z�՛q�o���L� �j��ܻ�~`ӕ&ͺ�v�@�_p��>�r��W��Z�T�>i`	%���.)�hwة�Uf2���=��
Xm�+���`����&�藢���
Gܭ]9��\�V�e(F��wB#=�j�8n��������5�,���
�m�|�Y��e�(�������a���IMA[��.[��VJ��:����j+NԹ}���f'a�i�y�����*@tNJ��>���UGX�1�  �.]�h�6a��Jd$�cs_y/M�_���.��0_k�Qߎ�K�v5P�s]�.:|�fD���.ͬ���& Qm�B��7��x���c?�m}Z�;o{в�*�3=�~�.1�l�m�_P$����y;{t�q��dy�^�NhB��t�����dG��4K�J��PO��Yd�n��4����ʢ]�|	�;�Y0brq$�@�*�z<ԣ�1����2����VrZ���(��A�W��70�w�h�v6�|Ѝev��	����=��oBǜe�L�C���o �U���-�z���զz��ñ� �+��+�O��IDj,ٶYs����]׃6_�|�XͿT�嘝"�Z�EE�GehV�[�ߍ���)%y��릾!WiL�z�*S%*v1��%����Q��#s�z�#�7\Et���}�Ƞ�#��mCFQt��
vz�!G$BN8BK�˼��E��;-���H���cgkv��a�p�1���Q����x(EG�����; �_7����P��V_F �:JH�[��5Gh����~5h �&�Bh�h5b�M/km�]m.��eO��Kkț&d��Շٌ�D��&�@��k���X��g��M)��K��w�f�Q@�t����~��Ą��}��}��z�ɷ���2�ᑆ�;��.�K(�C��*����7z�l'`0$q�u�=���uC�����U��1��A(����l:h׹�3�\J��9��+�@��֫�A��H�d3��pP��m�n�R�8!;=��ѽ17�>��}#B-ȷ4�ww��Iy(��:���q����K�͔�=�rW��Fxyi�f;a��j���v"#��7nS~
�S��u��<<Kt�*x\_�@�z��kv.�z�l��R�'�#�1(��	*R��$�W�]��F<ў�K���!`8.R�g%�xBڙ W�9L�	?�5�dZ6����Sڧl�^j�]�H��=��H��3�����5��n��l��Ժ�W��ak$���ω����^8\����cs�U��ϳ��]A�v���DK�{47#n�����M<�[g�]�1f����#�"��զ����9�/�MP�^W��<9|r��y���w8��E����S]��xK- KA�:E\�h�N~>��)#�� ��E.����$ԣ�U�,�[g�Ap�䶧{9I-���NΠϟ�AZ�$m)��_J�ؑ� �#���7�c�o���{���N�ҳ����%��Gft.m�ߠc�qgq(��5���|�����sN?wL9h�؂�SQEb�˛��XY�����}�_�G�QC�^�r��)�2�� �X���Σ��f�-;]@�Y#y#�US��a�-��:Ab��ʰ͌W/'��H?N�jV��V���,���Q�������d�)3f�����v��~ ��+4����������Z���������J�`T%��6۸��*�ZK�ЎC�PЧ�k�c�I�:?�������6#m�G�1KV���0Uϰ}ė�Q�կf���KGz����#;3��q4YNP�pU%��;�0o�k9���J���I}�wn�BN�F��M�	<0�Y;��7}���U�k���1$-b��4�S2��ӣM�DyR��:�BP<6%'t�PD�ιP2N�?�0���rm��pI�I�����ҵT���\Đ|�@N/"HU�&{�%[���@�u��%����x
c$-5�,��!��e&��`s�PT�����o���2ۋ0��,��w�]A~;�!j9���/ �XE��U�.�A�ʻ靼+�źW��_.	#3������%����s٘Ep�J�D��њ� �@�B$�E���XF��S��lڏ��N	uk�?L��4k�����j?e�Gz�w��}�S[ei��zM��l��]�����C���V�}�F��J�-c�3ؕ��M�c~�c��<\�_~�f6 F��7>�pϸkbhi)�L�ƫFUX[vѡ�_@<��5��@=#ɕ�k��_s��M՜�J�e�kH�8�a4�gQ�Y�
�� �OQ>y�
�Ϯ.g��^���C����6U9��?���xqdt�!	W�TG����֦ЀO�k��Z�o3U�x�u'Q��ma,�J-"'-۶��U"�O.i�z�p�C�/��\c���I��	t�/���
ԾA ��8��r�`��\���A��������웒g����YN����읗"�)�s�>�s���2����Jpۀ�&��_Wy�����z�8�j/�	p.�~ؚK������a��q`U��dfe����=8�Y��j�� �,����R��