
module CIC_mux_probe (
	source,
	probe);	

	output	[0:0]	source;
	input	[15:0]	probe;
endmodule
