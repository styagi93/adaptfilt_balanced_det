// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fvehr8zOZGCDnfVHDkDZua1hGHb3eVd6DophwzZXkw/lwzH7AzYiyEuNpy6CzssP
1d8MJjXYLvoSMlf+mggfK1+i/V+eVA1aaN7ySgRWoJgW/Os+edcgxwEVshnGu8u5
szl3zG+RjdUuLPvAQ/s/g5cF9rJUrjE91hA8ZQSqQ0E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2080)
s/uysFt5fOuyAgqKkv/vT8+nHkyDyN4bAnneSzizYP2XFEnj9bVfhiXwpZsj9y/g
RRHAJzqA2pBskhbIXV9lyIhIiUUAJXiv9H6WAwiSH6ACcSGy57H8d3lqstnHt4ro
mCD9pgGZ2bJdPrWBfLfpa5e3xT2JmQeLm6XwZQX5FZx/8c7GMV9C+lfcXt9+puYB
wa+dlYzK2bD560PDSEMq1B6as00gJ0T0iqLVbRg+PMeH/rOxGsyhInp++J9mRd49
O0yQoJjfP9aAYq/kAHjK3owHRpmnY2NnlJwJQJ9cL26ysh41dV6nILBf2pZwQPuO
/3I7Ve6bGBophUpWkYzIdiOPfroy02zzKfbNZQS1fDECrRl0byCDTOvp9sAys4s/
bRyh8uuSHgOM52a1GXE4+42bZ+XqOW6m+1t21bXb/rhlUzCeBQ/oleN41LT86Qka
sdFwjahe3vJYCU0VZAxGQfkftLPA+7KLAVSHa7kFKRAk1Ifyid5/yNXdWQcjYuSR
hKIAoc40m7IurHk5d/mH6oEdB0poYWtRm5zGisNq8ccyilNQWOR5mBh2n1bMrbrc
gbyiQ20Pcj6DDEgnHx+CIg5Jv9gEaxCMQVLc2YKy0GW+QkaCKvelIkVZrjtdPG7E
ASZQPxA1kdYZja1n9C5zfDDsJvNWDOzcZgWjmFXKgULUSiMllC3sX3P+/VdEA7aM
Gq3ddUMJ7cTlyFW2GNYOc7obHN04N8XfhL30PK994i6G7jpQQcVyHLW3ABe+CHhR
Z229kP70ATJh4U9vaKLm8ewgkD81jDtSLoyJWSUhXduEx8hZIXFxcUWO7KD7DO7O
ugLW8z+IF4nXUhFBk17a3Ow+GUUdZHqDLzdhZOsWaJj4wcAESaNoN8bRSm4HwK9r
qYWMPVBb0dbPNIAf5X9InHfrTVUCAwyUVwhyNE6CPHefT2TftXJdeyda1P7YxU5T
ZZb110QblJLjrY+CD+YZjT21jeulLmD7vEe3SwiPRLZn64efCWkLKKK/sV6Yv4Mr
B/pqo/a71lkLoK6km3jZ/qz1f80D0/tLYuU7OtPhdxXnR7hG88fiiiNPUygWIE5R
Tr8gfhCU9LGUfykqSQhkmayNrp9z5yddHhs58NPjplwknjutgRA5oMV59VahZafF
WiwW4MM6RDxAzyHBfz0uXn6aimRt2M4Rss4y8xVAH/g9RrA5yJswygXi8C7HEoOO
mSxhxLQLi0Hxwpmvm+pj//InJICpiZoYn3x2+5Ac0n44CupziURo/5RO5xyqL2By
nJgy+PslfEdtqSnrglnZyFTZ8YHC/TZNzeFDxv0/Qw+qcRHWLS+spGtYR1hPs0oe
ff4QDTipoARqQ9SGs+nfPereW1IMDHZL7tkZM7faxLE3AdBeMBQfaX3j/hOA0uXb
dVqmfk3MTGbkM6/jZwoLPcikIoJVXNmKXNoe+KMkn/7Sd4LJELMv08gpu25ID+c+
OYNFDYncd52fYdSI1pLdlhuwQFQ318M95eEAZStSvUR8dCTs6IbtYCopz6LW+1on
axH2WHI8yVrfwYOn+975SbGeN87cCCpZfKK/pWHsnJoRFUjYd3Yf2VBzyKzWXFZJ
mClluz90hvBdOtM/IyLFAidspO/U5Un3OWBzfYIVN6NMNEGUAQ/wJ8tnZ6A3PidN
R7iqZakgkoBn0AghvMmkQsDttHhf63gIqmaVnI+71FDFg915NRS7+50jQleIUrmW
2BeVce7d4Zm9nN0JW6hM2MP2O8TrOQskw0JM/rvbayRiLJv1COkT7P3OAChi05tH
A7vLv+6GGGmZ9MgztOTThZeTBWHgLNmZnKSWKKC+L000Wr+z8TPmrU321rYz3pr3
U/sxQgBlF9WEIla7Dvcnzq3FaOyK2mdu5MCRkxO7mxPisM6+JcBeSg3U1m5maYKF
xlxqMBGrn8mg3ukClSTBRs7um585sy25cubjViNYeRM8r4b6khJ4+6emE3JP7Q4F
8VGbuBuiQbZOHmqEwRtZ6UrrOYFBYfmN9KKzqs+I0UUSltqYeVQcexWUJQECCh8W
0Wbjr1geySkDKFxyKhBr8pHEdd3WJMBfDejQoc1pJf9bTO3hVRwjYjeVvzb7noVw
3SVSVNhADuT+JG5dr6/txgC11jAxiFLI3n2gAM70r2EafF9fnRhhN1tfXAySKmFe
v3rs8CsYc9TtEzjPGSE4hrShZKdl35x0ZXohzYrPmIom8QzlTi+ScjbVGToa2Vqe
qnWmS0hv1A4s9sEzsaCymhKSvnmFtlySJ3yPbm9Gec9qSvuGeXWz5/tLC4OH2OqV
w+veaDUvvQ9RsVUmQp6m+t6na7XeRjAH1GML/3woKCa1LQ7jXN5Q67IJUetZIwEO
IBM9a+QtqsZ48bsERb9Kbe5n6uU0ud4Cg7pkGODQ39K14/kAd7QxEidgU1Obxobc
wBnxOH2i/yf0h5OL8UpqX8RaaDnmShGOfDxq2l3VohVwu7NsJ/mbbCdA3X5DHKxV
MrwrK5AxEaWdDcXwtc4O/7u0WOWusciW+QFYjAohIiAByRih2kcPUwfL/buqlOjC
o9HBRnWccleo+W6pfrXIoHZoINuSAQlGLgEbBJn5NQg+KBg6auIPQ+GHoOQwPyoN
+lsMbIYzTCMAzLbPJm+vfMyNH1StXSBoAy61YvQ35skUqWb3e4TQxKrTVp8JEdVv
LF38ObdPy/4R8RJfr5M8CTvmKuGAipW8OBa6ll5E1hzX5V/h8VcURuAEdtolL1Ag
x4TNZjXgYi07lB+2FoyxJA==
`pragma protect end_protected
