-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sdONjldBCmM7YfpLvMMdZKsgec8DoF5codDWrbesfvBwCG0flaR8XCppLKq4UsR45h4KScKXFGWT
S+X3sv2SfSOxcd3RmcYIGa7tCyP9+a7KbjcIl6Fj9t5fF16A4nihr9p0387OOCkWZ6kXt6CvFxsM
i9TqCT+T0a0cevU+Kg0ye1lEfouWDD0gufNRgCSQKdT2RIOXuuYQMwukBC8Dt5hp9spnVTKyUdMu
LYLMr8YanBERkEjERlU2uVEn7DEtXh3VRmMPn4qqPWr/Ein23Exlz6e1ztVGeAqQNnS11Rwl5gJk
2FzEE2xYnErOKMxCtQhLJ7G4nggTfHxtpCdTDA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5344)
`protect data_block
o11raqn2CPbTAPqpb9MSXDIlndXls5zJpUgWgUenFBRyY3Y9tK0e+njfQhMGC0ImZUiJcBxvhfGJ
Hlr6WSXRXTTB7GpDuWw9tP12Efh/2PB6eJKH/EL0L4qOESX2WhwXoOkYtdVLwwHV6KcAeewMLpE7
Rj+3Su+EVxyKwXxaF7zVM6T2WKGW5bRf5AeVXAYOUSdin8ldQfelmasghNptLjVthYIgSGKUclel
cP6a3fcdV6jMaqbR19jbmPSH6rGZW5YHQa+dt+HunNzFvSikxqJA0AR6+2PMMAFnSkJeJn27sGwn
qZedRi3hqjWQhuMCiLjU6ZQmQmJZZZXCkMvEFJinaZ1e5iTqkGUiFolyLNBbMME+J3i47s0DpvFS
GyKUnH8z1zlYe+jwu+Zm/e4JqfWRHW56HmdHs+KHB792tf2vac8SHvECZKcUP2iLVR/qDqzOBsZi
JdCIsdzvrPH4Fsbn1tSIAhWh9fA/zAUMaeLmyA+Fm9KytCwNe4lcr1Z+4h03TUqbFwrt51m1gkWZ
0NvjfiP4ltIDgUVWSrrjfW9rQgM9MP3buejwMJ15Sk1Ii9A9qj37ZRboxgAzeiRBgaNAjRRzxKBf
fD5o50K3UUqrX4cwaAiKcLTgRIiz3qN8RXzDBQDO6KjWGvMOXrSn6pjvWUvNVkL8rfODEWMmX1YN
IqQnN9t3T8jPOU3QGkARa7Am4+JmtLtH92c6+59sWbGlhEvhIhYEkKlvIDLIJGSfF3V4UzhR1UeT
ZM67eNu8/lgh0Fk6IadxjvuWiq4ntSvuFiUQzsIvNGcgVKcmTG7Tj8lRNdi83H61g4d5u6IAHNfe
ERJitJA/QqE1gsIwH33bzXLQ2tilXVzzW4C3VXxQUumy/XKAGAIXZg5rBT910aJMf6c7I6pND3uL
7JYz5AIbKy1XbAtJ9p4ChMH4cDfnDEWc/GTeHNvMAxw0/OxXDmPeMAS6xRqJ8s4CYyKmhEIkr4XH
cUKTLQMMVXshpe2jrfrD4U4o+To8o40vuI6Y3IemZhbWJkQ+B1/KspyZQBWFeVZCkqbsmFb8z5oq
6QSDi7wfvNUQR+UV2lvp3rAGNrBSP+RCYx41WQgpnb3RixZ1azK3E7YD0CMzqVGk1EId8a2fPoOp
YfkptM2w1+M1cUTh9T5+bc9ThhJ8cE1WqSdj0Xb9WZU7NXUu4LfTqjgVGJUyKEcuVNPtGoviVpNB
XvvwyKttOUDGKPasmZstJEG1ASOI+jw20rwQjvg88jGY1oqeHAgjGAImgFcL0rmj6oJBq0TTOMvT
0Ni3ZjA9LG9i6xikqOs6LUa0zxhY1UsVOifKZ8w7NFw+c+BhtdF2Lt+6E6bzMh9xDnfe4EXhK2PL
Ubu4cxtqjY/ffjBTc15xK8tBzjdSDpdnn6S98oiVjSzuISvDr+AJMG4lhqSp2hWD/ZLcYar/Gi83
9V6nklggvyjsPfgivSUvSZrN9wv1EvIsvlqlWHr7VcsTLxF8ORpbbMFTtEzn//6tA+De28iM3Hnj
kzOLNy7XLIcId2PRhRc8L25BYqxjxbWcFa19uylk4Uj6WzcHZYhFZHRvFDtzBQkblZH6dxBNuIZ1
jHuchTvP5bNqj4LwcJ8uqUOMGK22K+lmQF+FjmFWAtlaCq94pSdazgK9Rz0yfaJGB4skShlXveqs
s+R+uQnTWVh14TZ7KDCyRIdWSpuFTnmsTTDl+ElzHF3Ur+xEC48rGNGKxKRibcND+9oBn4lBTY7O
otGJLlgaRsaI8PZpLoVuBZB2yxSzrboWuILwqGLUncdS5AMV8YxHUDO2OkwA7eeT2CRYvuSHUa9L
zr8LPcGN6YjUVtbWoR2py6KhF4pGZKpjeKLosUgbvv4Iq9rApL685zKvEM14qrfa+Rng//FMkIc+
o2EQJyDBL55CEY824L6+V/nMFZFcKM0X+K3Cc5Vu6+dTBXUUX86cq8VlPM9LkbHzFXSl7Pfjc3LL
yU1CTDAgWQ5FLpq8lJq9ug3JV8TjWqn/gmzGAsCQomHXgqoWJcsvPHokKNfyorJk8kj5screiz6u
oVjLXwDuPavc+G0vE2IVLUO4EOLtZ0R3FZVzFg0R/yHc5olZPwh20WTkcAbPoivxe5JpSjvm9x8O
JblXyndeaEkOZaIkVxMTny3X/p7qnutkSj9KeudqD19dkEPoT5KKXl8o15MVPk4Ir2KJnqBntb1a
soAJ+vLUp23Dq6TFabBUjf17AxS88EWWXUQzvmmqUOwXZpcHe68Rd5oHXfjrWPkcUn4/eluwW9wy
3aM+He4pbWY2CA7+6OQHG+vHbxU0HHe4Gsqe10VD20+qRImCpmJSkSGITg4LFj2TSkqZFAp5h/UX
nH0oCjqDXxKcpZREIzmHFQuDF+5raC/f4pmhc7PnJwS8aO5YXo7je21NrMbgZ3WHGxc4GFIu+NmR
mPjloy28lok7a1xoeWyXWjEP3OdGmWqlrCDINV3IsKuqUB2cd9o7uYGIoWV7MW8mSNai7SHVVsYk
V7cnVYes9qgoF7W4XL1vcocqYyCqacLHZOIGM4VJHDSNOXqDT4ZuzfHcc0fgtYBYrudkbjDI6MPV
9tyJn/wYQ3ZVADZIxrUlaNkta3GV1BQLDzylXZALyvZjBaXScwktVjuRn2zqk3qLvkMJuEvaBVrj
cneabhBSVBe5kISsQhvBsqGSF0RFroIsvLrtNSThTEOcBHUIWNTUVPytRySVZKXuxfnXEaaogn6s
1s03hPsqTtZGUf1Jnc175SXuPWSrCEf7JSl/xxkMHnokIUuJ3ySGZvqSu8bM6qaMxdifxNghhpi5
tPVB1tI5bsOxTexS3XyomV9/71OtfFtOw42k9eY/7wFjONwYVuc9QYgpoEKHRSlPNtgqBcJQG8e1
fK1doWVuso8E5YMWyJXNYrF0xDQDM7VRo5q5pdy1L7KQFsTFxSmUcIw1R+40rAa34JDJv9grxEPR
N9YpXGjVwOMhN9/MCiaJR0ICpiPsDkGMNoBYrihgXkRGjJAXoZlfUv4Vff9LNfRkoNqZHgsg8QJW
qMCN2L4h8RvKIMF8o52fGOF93mGAPGYA5XuTmedzJ12ScKEzaybBJMT0Zm9vUIrkvnxh5hQNqudV
qFMSVD+3Owu5huRLut5kdOqWK2HpgEg3l1RhP7TGc3KDVAmuf4iKW+qDVzBhKrBcO+C7GUtOiBqv
Cb/8JFQZJ0O1cImaycXYmsu5w13ruLQEad8FceOhSTXCACJ+a452jtzfePNiIVM5407VI78EW+di
7Wdekocvi6XRFGdaJydJBqGZXhJnnCUnXfaqpHhqwAUQ0nUz/gLexeaNpmF5lF0yuBA/EO0kZjSo
mvipccfWAw9FJENnJJN+ONwEon3iwlVSSbOJ/i07BvPmcugnrGyvEU+OutkcVLvoep3ls62bqMP1
tk7q7KJ5Q4zWcdF1Zop6jIeJ7uawoniDPNyGceRB5Fal+/zhjf7nuzN1eE7GEuANwxf3P3RuYD8+
e1ZzofLWkOgxp4D6ily1G4KsI60K/ytP0uivznQz7jOYiC1Lh7AvBHT8MJghxv3oUdx4pVlRugkG
QVY3w/9jx7JyAgBjQ6fKJiaLKWf4wynpZovWfvjDq540mHZ//ngdGMA/aAvNp1YNKw+z35VegG2f
+i+abmJAyLrK4lCsKe5tF3Xeemf8ZbjFGQR24yGPScK7TicsiLc6RDSRzE4FJnnZ2J3dxD8kjdvT
Bltn57fQTYki1zgWCPAmuPNRrQkajvaBrRc0VXYQ69sRFnot/pXIIzG5TfZWt7Cm9DNxz2W5mmoD
523K7zCfJwsiH8zi9rSx2RW/aqr0XP8aaNaHCZLDnnuWY3Qg2EoFkvklyQea7RMp66CvI1SEldsh
Fi/P5S+dhUUgCQRas3Qo7kjjb1Sv3nDh3QvDJVmuiQxZ0BJw4DHnLarAOm0UgBIYPgbXSxZy0Ss8
nAmvY0rgIVPsr8gqM31gau/wd3idEBrLaxYJFklLjeKrOEb6fFRwSuq42u4E8tklPXnOXKnevjGy
z9vouACDbS96B8yN2MNGXGNPKoQ+A2gqtuQ+rHd/XU5WMFx3yfeHbtpB2EtFgN/lJJbt8+4029du
h8COVICHRRhgcco6jbBDuzbjwUvzg9ZcpgUiMBMSGv4tJKkZDrf5IfMtDWxWkWdNf6B71ty/erom
rcCKv8lyYFqlrUupuOGnpJGexGpgWrgS4O9BayU1vrINx+zatNX9g3q0xKYccjGB1XrBWfCuBp/d
Y8IwbbTvs0YAU5WxB6BgunJsCTwwOhZ6jasqw8KJ7UinyQ12wlPBGO2zCP9NW0aaok2jdG8JyLRg
yb1/rr0iDzV0nlyjllYbihXQg4D2Zl5fHakIzOL/QWRMXRR7D65Src9BnN3bhNb6CUV3rusEXn1j
ImL3+PRGARIgfaT7cZxgj3yOBp5YEiXeQPj3+aM+/fEWPju+GxECL7InwLNVzVnPMWHvkCtJSbCx
QyTBASH3ElXjWD6aD3WqpGIh3yHqkDG0bX6V0OxNMZBSz/IXV/GUKJc1nDwVS0zHF7aiqT/cS0dj
u87p4YB88MygybUeGpa+EzLi5MzJCxgaAwN6jzVv251TYmeF+rioCMRahXht024BsPhIssboCNY8
8rM1/TOJ7q3ZzWVgqYBeEldKLr8rAsr4qyosp3MUJVOJoaILTWXuwW1mK3p0xqrX7hSFawpJR8+d
Izv8pHIeRZ90Nuhjtmh87uTaIM3KiARxaLoJTqXtbBbfhuHOUBy4dYjkuky2PORxK9yrqTPG08ND
5pVb4r1kvYuMA1DVbignMIjsRHs3t36QlRGIUxCx8/QIgkmQs3Xr6tPAQ216tzBtCbGCatXxClC4
qoemoUvW0Dx0ra3EJCOkD/CkAOp7NoPTHd3HNqH6m5g3wjYN2RvegcU1rYVKCOfoBPJyyOFhbJPQ
ZFZBOCt8VG99MLYGqEWre+uBk9mwOHgw5Wm21uOBDWDwacXBktoz/fntutwzswmag0DsOZ58bhel
61eaIHvhNk6GArfpbjp30llPhh4Cu8c+dKwWZh4ldT5d29bibgYZyMFDMa9AMCeEZwYTEtXAH/4i
Lm9jTlw+x6ozXk4eszBiHFu+egn8nnsMYIGJ82cK5ZpEFYXPiWvrnMTSnC1QrLjt1H01TUBu3oUz
Tn1JSsO8uOjbiOTR4wK/2mwjyn+/Uf+LICi7wy4kXvDXs5N0gwHHcFFnTxI6YmWnG9o4EF/9S13Z
8Iv0nGmaJG3jv/Ab8jmiHG8IM0Try5xKwhVM2Y2aA4UZgMERvNGKL8N32aVb105gHYxo3jFj+cdX
XyfCgChk/2v3tE2sNrROBBmAzYe5G9jLBo1dfNrsmGYcFOtdN0Q/OOe+c8EUC8aVbIWzrEGs8gRh
XyibR4iCHfec6cRnXVna49z9YhHa7swPK65hKr+O1TsQsJFQF/rTsrUL2b+Y8q17GgAh6tA+fgnI
9nNRAuNRpGTtibtTOkGLeZdr2Ml4TAn9XLupHsSouej/UUXQKsJKHNKJ49lmCSovNSJPuJzXR5sx
GRxELUlct1NgRUSdTVtPbuWY4EjbMbVE1LqEhdbfQ86FpW/332RCcFeUHqbE68gNc2KZ/EVJsyih
gmpTNCsPzsJBC6Qy3z1tQyoMAhns7XO7G2lb8vMHVSQwLGHFLFYa7COXAY0ZvpiNAfD1mcCvZfRv
L3R3s0MmzFRZ68CJhkfRKjShUsiswhquhCyzYhmd8a/JWStuXVqZx/9sopyXch4Zld5pR4GEugLJ
rIsUtPunJiRywuNnkvXrWbVuCGkbmkvSk/XDMA1OdHtn1xdb87W8oTO9ROD+On83+mx91uNTt8fh
kdFpzQDNrDrGcJGcH4darML2kBbvzTDfzOfoqmq1d6p1+dbeyA4WkeRof4JRf2VFrgGB9CMozuAK
2+mQz9vJAF8KEGkASbtAHTHzcJpXkmREfrs0gbtu+BcxzGqMJ9GZUBP2BM1cJMHoYgNCFVASYtV0
ArRtF4eXdeqH+Z6sBlDfxc5eDu56myZ4za93gizvqn+jAYaip/U6HQEyyskR1hMEQn5CA+oPGtoK
R3+YCNB+vDfPx/zCGQ6GtJY8ggp0F09Z9sdYdoh26sKfdFXsXyP5Vs75SYuoRyHk+c1xxNC7zB1s
ycBHBLjVCTNfbwiJJSt56YLDuWUVzE4UYIKlwQ1nMZZ/1Qu23GARuVHKBTkHFcFQa7U9aTpUQLug
huMkXJlBe8OLRYfNzPPTgTgHhqFbWxxHzyPiSVolqe+sH0Znyqjd96VjfHxD7Z0m075uoK6lzhv+
EPmRd0abVeO9b7jpJz5KxCihEDMSq4/fzAYA6AOiAhZ2ZiRGtuQDhxFhfF+TzPDTUgfJ599/4COC
y8DhTqwrR4G5fe9d11ObM5cO+y1B6Tg9VXVAJMGLpjTkWCkbj13qfk5gcr1Llt8jjejDQZmIk9qi
IxWahu5Qv97UalGW2u2c6X+ACi1zpg7BI4jLckziSOwTlYrxcJILnm7CdpFoztbPbc2Xoc6JMws1
xVX564FI50mK8BGu3eotIvr5JOMY8knioQUfC17wjBgUTl7iHjakNlme0Lom/QGNE/zqGrtJDRSN
Rvs5uDxsttNxGvfuxP6/UTjBqT2M3SqocXkh+JCFPcqf/8NfOyXUO4wW3ycmPUUS53W4E05Qwk9f
gJHjY6hxKw1XX1v+6GY4yzMl5d3iBgsuGpjfdRXetAQuVGEr42E7QTH2JjMjMaClB6rED/5dtrpb
D/MLhnQstlBzxe9lhWjVLfMX1Cs4SUn77Z3OuuYh/liCUcB+rzEWwbuZlOOvPLWshQSx74um29oL
lHBoleV/tmXVdLp7Re3sW0jvBs+7vonGykGQCPo1EKsxueq4q5tERvdTbf9evHmE6MJKJUhrG0ur
iIH9N32Y1R5DxyZI49JtpKLbCIDWrvzsjmCecYFuM2MF0UvPkLCqtS0LWWNRFEkjDJ0dohEUqpGc
G+u4P6enfLuSzHomapafghYmZsssBGhYfjO/8tQFpvKoDPx3Z7JvBPuJCwbvXeobvZqo80BcwycP
W3Fxk159m+cunlAiYFmkPcj1Vv6x4U2SlX0qrxQnTEhs4ZKv2BQVvEvWaw==
`protect end_protected
