-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
C+tGr4ZuI1bhLVn5KYefRH7wGedl81beCjVTJvJNzNDuHhKKEtqP3otGXEgMe6pO5Pu8r3KA8u7F
KVqJu3DwYme0XbbZKw/NH+JDyTm+K+1UOOhu21+V2Iok3BmtOBbK6+zqydCyQai/szmZWe+xk+Vs
RQtp//XFSrNWTZui8TUfZiQ/JRzSjwiqRKerrF5+7vVIlYnvtYrTseYTio1WvQfBU2gY3siZnRPl
Z4ipLexctT2CmqWhzIKHKkjYG33sMUekvCMFdjP2KeLDRikS1n8MsPUafztYoepqKdfszZf8B7t6
KuVqUUGh8qC9axPOZJgL7oNTEvytUCCAzpqaMA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
wlBlGXf5kYSFqCROsHj7xfByQ4VII22fZQsFMU51lGmiOygg92F96RVxMoefLSYz405DEvCeePni
ScF8Rf6DwwHCA67P0/iAhkf/ypSl37j99lWmvpKgdq/ia+ZDLXiyfw+jcgp3zu3lifzdviIpEcgF
9EMYQyX09Jy1+frU0Fr5k/futBKoFHpGXvw2MVKMewy1oLeYRZSBAO9QlbN8r4JJZSipL+cyAkjs
HGyLoo0wSnNMZPPQ8WiSbuwIdFq/+gk6Gfi/hqQfYoY7yt1Oru6xtGL7HFvuhRawZ0CgCqVIeT2h
h29ek/2OsonKgKmnRd892ooDih+lM6MV+gs+ByyznecUC0vnbngABX5gybgT9ej65cpWvcUH2rcy
PvBbQULFpZNUVJA2drbpBgzaskCRmDl8xBvwS86evGXKm+ug1sD8jxY4nJAR5lvkfHq9TC5A+vs7
4WULFADb7E/s/nsYE4Ijt45wIW5I/iqGEkCqtz8v1Tb+hPclLowUV/05leuVyZQN/FT+fkrqyUBk
PNFjN80tbkUzaPkDVomNzlDjj/o2pPBGUZy/9zjpBQeVYF/5pll+vH1am0tu9PP300N9SLHRjtWj
KNIoudwRW3GIYTrf2cjOaFrK7Uvsr4/3y7VLAjJLJos0bniubDB3vGWk5JFgMsjopfBWXrVcIf8W
3gQg+tV0BqwWlfIYl+6fDLOPMABMjnrIYsDxYU8+bFjl17KkwJKz7al6GFysqwbqSXH+aKJ/eE1T
Xd1lxn1ILjF8Eyr5qQ7r3w7vymegFDUusdY/t1rNCWrdhjgGa9PWibMEC+yiEij3v1R8mAIq52Tw
KzJNW+kLEPF5XdO44Y26BbsTkIY/Xkf5sDY4DIClZuls+h2ZNWhLrJsu5t4siBTj+FQAMvJmOUnY
PqhRwHIxgwcolLbgQjWVTyf/fJslDulEW2bEwle/GVdVL3AJ+/NdfiaFvWZQZvdBJ2ZODWGnEkXb
jhSAgk4FTiA0hYcqwGhZgAzqMCv611CpNUoIyKwOLMyZ0e5ks2+1JtYgGsif3yP/JRVFNn2sONue
M8ztDHJBNuyxfxtgVYGCXXOQRfzb4lH+33WQuuoeQwxRCNAGyybBeqgzd+UtqVNN4wnJ0MAf49Dk
ISmcoYDrUzUjkHzHA8y5EK4zdm5ZgF0vDDZYQKmYn35+BJHt/Yr1lxDEhUynKmHOHhXPNmS6iGfb
SH7qjTgPbpvZa3GeaWbBdPgnOBjhXsqMo8oCU2y5IVU74NYq7hHg9YCl451FzaBI4GYxLyTA+W2t
oIedL9oTsX1VvJisiWBBL5a8rYrkEZUTdfX+6tCiiKJLKUSm+fjal5Y/9ZXxb7GxxfUjx1FgcL0l
VA4Fox5Y9ECi36e1YhTWESEJxLYF+NAGYB3tIqnkyQAbXk4ntZ4e7ULVLgamAwj7z55/UWWxU51I
gHCikSq7h0YOOTdgEoWXWM9ZTGsKy0FKosnV3eBCfe1WLngmMYg9oOkZZTM/yCA56WNDTQCjxIeL
1YfeSVe7P9jYfQnAdbGeTQib0hn/3H+V/COTo+eXKzbbnXHCKxPTYNV2/x2wl4na9zjqy3dIBAXX
HY5CAcyb35ajsADlFkjWI1ogxG/fjQxskUezUXymN7EfZmpUUmUzbA0pw2gE7xG0kKRErrLz7xnO
L8R6uMyPqwhfl6uM+w9swO3F6n5BLu2dBVwsqPfHiG+RhRepf7GA4pyvNLxn1mB1YriuHUo+5OLf
3zRPhUB+EscTZhafe4WN8hVPLxdO2rFr0C6CkDmIaJvRw/wrjQ/QEmiF6J70gjWX2x4anZ1FPDEt
iKZbCmLn4Dq0sEHm0XwaHq1XYw7Lq3z6B8WMYfeAwNvZx0EFSYwwUYwv0iFiYq7Oyc4fSq9z+RK7
XEtwhdcTw/kdX1xCO5T5NeBz6fHdNzSUvRKPzuKh07EgEh5sIrxBhkD8eEuLeGDOt0feQUO2aIYF
5T5JWXdk+YAZX4tjEDSQizLdWcGwbEajhtWIxIj4CWRg7ZzuM3zxg9niTUL/xllwi3BdtD7n+7I/
MnnO0N61OcYC5bUpe8s9vrXILNDJu7s6tW5J+YVUC3iHs29v3FIRnieXZmKnYZU60pObPEmHT08Y
yEwK4HHUVoHtWvMI/NB0qJfkh6WQclS5TQZdGTvvwh0rCYHxTcXWNH7N2TGa/1lm6GT8lzqlpMyA
G1T3xTABiQ8c5vDBeFnZIsIOEFoLSO/20DFELa83y7EvwzPXBD2DyezMDKb8xpYbvMGGrgJK8bl2
/d73e2EU0UUUOmJ0x13r0G3b/I5EsT+rd+6y4S/JTedzIRlTt6QAoKQqyXfowMpUWAq9UvvUJOpH
0exB95b0V0gsvuxzVVPahO8Mt1jpgQS9QcIgvYoTEwxH6elESw+juIUsN1fnWRk4dvixRCKcv+s0
x1fqlKHfnEChz5bH7QYqlUy8eFRpDwBVh4sge58RGBO+JpahubhH/4ZuIaQjMkLd0E1SVK72PLcJ
b9tufkuPtbUZlZbJYUPGcWq9I1WfYrH+22NVWNZv98wItVdhFPSpJCgCNFtviDqAgZWbHimDziKZ
L12VWAd+AeH9ZF3+O9k0IdzJOxj7bEUEtghffh65bdcn5Og38J+pd6anObxpyz1JaSIpYUF8wOzw
6ZUzyAHyauZF71WAjyMrJm4hP27iStXPGpXE90KqLjUcuihQjr1TErx0f2OJLzC5PYJadKwGjLqs
Kv7en8Hjudbj495qMQIinIEqri3jnSad7mGTSpYCV2Ul4+lKPmFpuoK++d/pjE/lTs48QDS6xykh
R/LVq/YHgHGMvaHjHKUy74OcmF9/IBisFMXH9xUGNLl6sU0/VWEUpqgkwPiQIscZhWIYHWype2Z1
0aI/fwVDxFseL6kjfm+3GTWJpYQswUwq3+0NtVBht5YbdwLFqKomSkCtzBor9/Eh2w/3z7X77vS5
2gCpFGhJb8MZJfubWMNM1TDui4oDgBGB2W84K/D6sI85M1JoXOMJ+DYcuMUoNPMrVfNQYYL/rcEl
BII1HVYj9R77HMqm/9buXeY9U0oEBylcUXAii4Sc4RMedeYT5rMfBsbGWEalBLIOfIZEpAtsMhbd
xfGb+uArLL7ioUSIb9i4GWtrLh7w3/qqo1ipDVRc/kxI4l22eFkATSrGekhHdoFCIRXHJmT/Cu5A
S/RrUMFe9cVwjinW3A6QSQocQe0o6+5jE9NYmk8aKWp0fSMDgWDbPvL/THXZgt13GytA1Polzq9i
bxwrzBCrQka8HKpG/EsbmFUGDVu4ys76at087bMAqCbkpZjNvLQqRIEy6Y9haEH2sACQNijn95u7
VSaipXO4WZd1z/KqguwnSjjLqbMTyX5t2+1DTOUNm1+EzVEQ6H27b7/7aDXk0OuoNdDjI45euBfL
9AWylMZSbxmHxM3xkeG7FKCHPxGg2sSWE4UTXgKGbYx5sf9iTwDkW9c3LO9N1r/8RmXfWQAiB3iK
FRb44+m6VDYSZtKEXditY6UUppRYRZX23AS7gjzwAEHOvy6KDhR92MtJof4uRyAI0Vyxbipplqcf
xnrSCY7uMPA7W4DvrKqPNfDgwP8iDQ6ZD6a/0GRY0fNeA31r923/Vzv/ZdhSHtlVXkJoFxcmvWg2
5hItaDMP/afVFjNNPzqgIvna8f1s5hBiTdXn9MqzKDMbhkh4gi9SZhgXJv1MFQmSST8/AldhRU23
xBmukA5DnqNHOJZ9SfRMpG9l4CCLge2aFjmVG/SaJd3jc0vnaq3HMzsnkb+M3lG4TCM6KJ+WpiZv
XgvodNb23+Gsj7/wexe5q6lv40RQ+LPG68OSx+eTY3q9b4/H2/SqwGnEDEZ1NEV586DBWiPuYcqd
wGCeJBREsacSI6yznDOP/PqbSde2j1XC//qCyoviUPDsyzQCLHH8dMOojG6tc2UxXP1J3UdYT/39
PekJT5tTdoxd2eU8E8G4jIiYvYaeRjNewJkRsZaREq+nHZx/Co34ioYbUH99PkXFme1JvxOqCXvV
zxe3fgg6wX15fFWGZLc3T9CFihzvjF/A/bcJ6IBDVUsgD/mgTpfo6YarBPIgVjYcjDvDJK8YauWG
fWrkzg4PbdMIIHqMTpwsL29fJzj2kzAcwmH8QOsmxytQff+k78n2L6sCg9wacboAx8AXaP2y1FzA
Di6HRxwuANdCqfQbJypv0dGzDkMV+D5N3WcrmbkaazYyihkJnXbr5otBh1uphIIjhexF15CpSP70
4fS/zffqo8ro6FQtp9PbphivIqyMH0KdNNEZLug2fGG0mKSosVHKOsGcvq/1JeLqKAj1vlpaz19Q
8pEPnN/YwGoy1Miegp5+HA15MRVbdvExVXki6ygEsAmJDPf3FMG2c7JRPAyWkS+fMByc1qXhpHkQ
gpZmCS9AmNuKRt/2Vl1GT5UGEmjd3fKR7HUzySV0kVZivXuA7/1YowEUe4BKUNth1rC2j5iGRp1Q
5flX2d50o0RC7YPzvV6GzdB9/sRun4KYOB+7Hw9vUSz4qZ5pnsvf5b1dHcLEm91OKgHI9CSVwjC6
SIAgcXS3qYRw89mInzhQGbkhMo6zs/vMps5IOaq3qaQI9TGpTqF0klGSsP9BVMxgIUcSQ5mboAUG
TuV+1qMNTJa61btJjFWg6PKWpsgYLdJXHkjQTa1uRHV7xA/U8J6Rp5voWa7Q4OK+Du+jlNxzHwH0
8BWKIsn2MzJjXHaXYg6ltzA9ZV7kF8c5psFU5Mv3KXCuUsfTiBpLRT9cPRWj+rrbrmtaSCQYF1KW
gMkQQICJfxBogBmu7QRKfxuMk+TBYOzvtp5188igAWM2VqlRKaWCGdlczpzMybd3PB4lkCXQf8CW
aE/TMaMfTaeD53aQ8N6JgXl80LbI/Vd7VY7v75KKG2cmpo+c1cGxC/J20skgWb/So1KBL4X5R14c
Kcb9W7CkB8Ptm6HqhJhWqN0BqsMmkisxK4DZz/mIAnxyrQczb6TZBju2bkoNKQisRbAz5g/ylYYg
/P7n+fcAPhk09/k2ZRX+vxdgU1wfPV5XD8I/djPzmk/DZfGgR/L4ZKHDxmU61Wvn1Wj3PpzNwhUI
F9T/4YKUQ/NbagHhcyCbXEX+Ky9cb3eKPHxu49WgYmjtNytomMnGLOpU1ysWrKS0cBP5kHu4ZfNH
rbtvLu3haUN8SgLGclk4jFKksRmx+opuxCMJCPi33UiqaxWPOoUCxCKXdCombtyknVbL1Bx19o+L
kAFvcfRSsgH9Rla17MBnjDxWQJ3p6XLVA6DpQV+YSa/O8jKtrjc3kp1gRealcs7TNZLWl9Abr7go
7D0bdZvtaJo7SdM3RypdBzmjrR3g/UtT/YXM9bWKSCe1BP1K5gNyizRZA8TW/Hq0tBmN8itLwR1N
1L5mtwnagKAuu6TARjxCh83V/TbKRp13zOaeoVeBU+Ic8g/BPmL2te4es9A59FciC+/goXvH91fV
yfzkLIzdPIUgD1woLaB+bdP4Djj1PMTv7bMCy5F4I9DB55+BUitESjfrcfb8F9gOcuetGyrWJ54l
mASv0ZrnFV0kav+q2/YHqDCFB8OaierAqbVZ3kwVcqqEz36eGN7O/J76nSEt7T0cx1NOFDPdHV9v
oiYVbONTt8YATV1QfVicYEIAPpIQef3g8iq4smqnzpW6hmH1TDCm46/G688ekc7Lm82KRv4DcUTN
5ps4o+/mTeTMF1yee2RVXpSuEZDtnEH8nxIvkH0aDOuM0AIxY0qjd5A/GoMZ5oL8HxzjMKzS3IUp
n8+2FyHBttHZD/DbeLeYSNAGbpneH3Rgk4d8vhwxD6V1k/xD/r4LrLziFlEuecShN0EfhXvystKc
oCgotWPzDTWErCNwXr1aji966XBy4Jv254mYHwgyelcXfCYSDZ2Pf2sdOk3/gpaz8TRvc46LrZEH
AoH4J3mceBmIF5dx5LUj+6JlbQKaUp9JZJ0Wm/yhxzDrBBhEZVcnR+Gut6ogbZi5pjq6r3Tqcl5i
Co+PV7/iAs1bxDNg5ui9G/69wWfUkZDnK/27dwKt3rljvvPrPJiLtnV+kvho4obm1+jhktqjWMHk
DR914tZzP3NHwWq4dnglfwy2i191xDZi4zoiL2022x2lReZDVCfTgFaAUUt9GOXAIzwfNcMFMJB8
VcYI7rRqcVgtn+Rc4eXSA6CanjnYG/ZWoc0S48+wJf5BcX6TrCTVMSbUs/8NjugySfP7geEswKzb
eHsIvN1W2r2BfWgIgGP2EieJ3srCcavzGGP5cqbLCHwWAswMTpEdSjCytYCWR8508if/HufkR20/
QMQfPT1CyhQWHcCvv3H2WTCe1MUZpRhS0D8UlAAcl9N8FVi7PtCc1WGuQr+7qA3hagTO44AzVaZJ
tX5CuKWugBjFa/aNlwNhXZlHfMrIQ7Gwf1zfdQWRCC83uGGVxjxbNLl/fSRBLsEMh/EI64TNWZDK
ZKRJWSb6ekjFeFKcNHOQjdEc23D+H15kCpJAO3z7MtJu5XzaB1htfiRl+zVAk17G1xHCszle3tD8
cy2kTCk1etKPbNDESYnVCwQtC+tGqwMSFC5oBmRyX60oPKNaTQhSybFeyh+64gwC/uw7MDHusmWj
dfI/XOELOxteyinkNv70CaSfArXd0DlIiWNLaqi1qs4+Zc7kc8mAXsGuWG7tmGsoIwGEjopF9eH2
1w5j8u4lAmrmiUFfOdLpN77tNsI9uGsH0kRytFEnHoeESBMiY3bG07HhG3YiUOKhAJyp3z22XPn1
OFaNmKU8gsMKmSEVdREF9BcU79uEIBYAhgJwMGdfMVyrKbwH6eNdwsjQOilqyKRGzwg56agFtVIM
QrYVslXFTlNR+Mtfo5As4QRypafYgOV9YsqLw/a9vsvKHB7Pk+CWggIc/wNW4LmNu0vp3OgjQ0Ny
EmM0SYNO1t70/GrTQOkj80Q79FCLeMsBeA85up6WPVquu+tbujcZeRZM1ZkHrWDlA4M+c5EdwYZc
Lu4SzXnnPpli2jeUnkq6dcSN+zDp4/nOwv6DJ5wxZPl35mTW
`protect end_protected
