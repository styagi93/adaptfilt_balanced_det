-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NKE5kvv7F8YNC9gz5Hq/lGrYlzid6/6tBvIV7skKfPFiJ41/uH1OUEVhBKwVijxRt3JI/T8N/SwN
vGOwc9VnRjlz6CO1Mc3nUGhrOX2sQpqwL1JRcp4dR88eyHXq6DU/oDiQFVM8gryNhlHc3z3qZKDH
1dgeAAFsU4eCtq9mER1nxnE5bML2MD9xw9GzsmBtjGJD9YaA9e1TfKtjQaZq0ZNI2ryKJQoZRbX1
W+gZYeclygOqvGeqqcDmU4kA4WODiZ6zwDZKjMFjWeNZHBVlFZIyI4IAxy8hhM3UCdKY1YwgzV7y
QRO1rkWtwqkvpSeUjU3aLxXt9GvSH1rIxMahkg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8576)
`protect data_block
gF/stXXSkV5dWd5RuGDMrdJiYLM55airD1K1TuMUj2K4zbfA0fJTTRS8OvnQsXqy/puJbSUorhG5
STrDCRpfZIHjnqCiterFpd6vmdv9jKBPT29MmuxTd5St4dzGoMXpIWNZfdzktB+hGveW17NpTeS0
v3x2Opjvz+aLeWPmT33wObXCG1d1uceBWJPiQi6oZu2P9QzsawR5M4ol1Cy5bbMfx19XrprsC2Lm
25rxm+EjZ/FgRWNqKty5OA092BHyNfegBL8MYbn+Am/K1GyzOP76uB0+zXmkAQjLo11QwuD8gZbx
+h/M8eKSRJbog3OdaO0Jch5vcuHwQHP0vRkp0Yko5JQwZoBy6fQMnyTQzVSuee09qg0YDm3M4kRn
Nrt482gcBmovJkOTD+OxM/2Po/7pVihbm/RnIbOQ6B3gBaGPc2BGeJkfGn9F6/NxHLGvMMNDq4Zg
EITAZutmxVQfwciuPcvP0h8bHj+axyqHn4SckIEqnsJ42nJe//H/R8/0ro7a58XfVbYNXhagZeZH
GvryFAguQUyn+DXfrctQCmMkv1F/+YNvNfG52Z2AJQWQ/IqX86UBAEJ2UM0PWcAoU437TTkF/gfq
80UIFgCETWHQgfEPBVAfNeLv6tCRGCliOgjMHCcaRoA9F46ooZ4+qcthSq3bG9tkGHPamT9VgPtm
ByAdAKJeVB+HHqT6jb0tbd7LpzB06QFUaWXag9QQzOFI+L88orQzvPYdqyJAVG1pn/NBzE6K9KD0
XHoNAeAOiFXdbdvfbouZ5wUpNnRvMK5Gg43bvoO7GNf/zh34nf13adshFQmzjghFhH52dRyBeUvd
kYAnAQxGNMyc7oiweJp/RWA1TC82VJSeaYrtNFhSbfDZ+KAQ8L+6cDPofNb+vC4mbMNBuGXCXkvN
KkRmtTQ0kk3aWul0KzkYRW1GQlm4cP3MNRajugTLKZGjX/2ovlljb7MVTrh3pvzQ7Vd2ce7kXxRM
aXHwyctYEsE/MqoY7AZ8aIQQRPkS37D3k8ROaJ0XX+ebBussAMv19vnlp3rQtKE9bD6lVXWu9V3z
WAUzwn3GM0qvg8EfiTdDU+uPiR52l+wpjiCPc1+FlbsJdktC9SjQM+ZBaFB+IpLyAm3YjuoGgVCT
NU3zYcjXVSkceTnvdDDAQualnJ1tsC1LdPsyzndf0Bugr8492cH2eNOEWa8RQIZG/IFIrRODn3Ev
V1c+iMfMBHlwIyi3EA4Qe3Kz1BCKIz0qdhZMXYcGZkB3wDmA6M8zD/NOyQWUoZUFdxQ9xaN9lymr
SSI1NzYlhaeMn5FbAe6AzCb+NjP+YgRpzWpAYsN7xSj1PNbVRMsJ1ecqekBOJchtuO6IXsl8d337
85+GqiE2QVEytVMNXNogtMtZSjSbCvagdnfw0sE1qa/08C0ktxz5Zhr1tBV0PpYGCGQfBIohADdO
r5VdzcLNlDKVUZfdUq2wzAgm7YLJ9kfHKaoOsav1xrOzunPVynYz6OyHie0WElE+Qp5c+Xpae0bm
2RsVgDNeeTYi0kpyNRoNmvnGShHx6Cpla9kTNTyBPwu8dFaOHmtZXq7iE5kyyRamWmZttihS0eGI
1P/3Oaed/+uQJpsUTK2V9QCorZsor1nsl4BtfzSv2ytoOAchdyVGTP3AFH4szzwLd1I+7ivO9YoV
fu7sdKJcEIebdZgM/rNl9Kp3A0O2XDW/CtGQMWnJ2vuJ1d8bY9hNyDmAV2GCT2WtS79yTmLU9RrN
F038vdLBWvALYIYe2RLmWWgmqn7qhKjp7g+tIzwIX/g0UTJLfTT4XMKf9Q5r5p05oTytyJumYL7y
DSLWOIpq2K2ztozWBLKgqmEEdu1jrowXi9NaMPc9MmgeXR+L3Q64IgHd20i1kDTBilwrpwPFQsMo
5VvSLQwNvwPodqbhmEpQgLAlaJ9Iy5e1AWu5v7LHGvlFod0ydXGlV3zemVnoXjOmYspouQcO4S+U
9wTqQK9lrLEYdM9RHvYXLkh9434LznaIwOEuibsJFkXiLJRxOzXtczen6QeH9EcDaCyfHHeG11RX
z0dcf/79vdluvVuNVGR04q5e5E0Jm8RpT6BwDdDrQbv2KH03o2oDFS4/xb5FgbomcH/AAdkJav9x
JUbkhBQBPX38G/pHumyLp1wL5oPntVGO21Zw/ZRgN35NDI8qlPT5Sr2mItjJRVYK0DDa66d1M7gQ
CiTjbaSPBLlJKxkwtdbJwCdiXDIy1o8hmsBwIiV9joiEaf9hwcNzeIzrjuvTWiagcjwtXn5e5NDw
WEVEMYSfjd14XAks98YqZX0oirqA4uPn8s9BM2d36wgbIrB5WiITJUaGtlr+JEO7icITzrb8JsCq
RCBp1JM0YEJmOwMsmPGNXApQaQ75zTdUrBbTpB6N/eUhhFgwdXeHDFffkmhkMr/8/W9DGGlgD7YO
VNtFMdrm9n9r+IXPR46ZBT0eOavhaIqivlTsPk6V3ObHs7teuGhJR6g5Cibfd6IgTyGAvHZd+ogV
lL8qlld31TQoc/rWLtI4q2O6l5Vtf+LWTJbGTOYGkADjxW6jNKaeUv9K5DY5Qe2+usHxE9uXhO0k
wACqGpt7xQtiBYmkcabxMnfctLZ334rqeNKEPgnhwVj1SEDwXuDKh8bjW7L1ZgIO4CWjz0K2SrW/
QoKOwnnnIgX7kS+jYAUj3aZSm9eOsEETXSIaNr/J7oHVtWCcJ/p3bcT067UfLBVfATL0SdhQax0J
w81ad6VpGaA1u2JxxIMJ8mce8IQekNYYDjVvdRbFoerjHvcZFMp+/4/SGlnY/hTnMEWGkmwwwpMD
f8g2LEM3ypazMxHPUCFjDmQFu9i2kDuTSkA0Ok1ikVmJkdlnOcKD6uGdux9nfEQMcvd2R8BW0qOe
PemaxYYGQt6Ys69adr60oJ+mWwJKg7u7brfNRwnAflHCwIV7hX2NG6Mi36LerjAxwN+a1gZA/GJN
MAGNM2qjQeflyHDZE/ZOV+WLK3GthVT932mr3BgNJYIYbN4KiT1Gzig0XbMeslc/dZXJA9FK+yuy
9fzvQhXmrAGy4Whyc818E10tOYS4Me6+lrEw/UHVVwp6NRFe0PuFQr5PmP4nG5DbAM8X93cOZpcy
Dgxuf8RkQs5s4ooFIN4nKXsKCuUWiWOialbz8x8b+0ZEnBDNAlvJN1rdAgFdCJW9atJM37dwOwUi
SSSmPi3iLjvlWBdaOa1rwHE76c8D8f9BASUv/FhoPnThGEXMUaAY06niX+1bPjUuUYT9BvGv8Who
LB0tSdHvEn807T6LpOGz35RRKtPFQsEdZP9TPsPG4mi9vbvnKm44kb+GpNmviewsKG+jxb1BBHzj
InIh2tm/VB3K6mUtzFsA0m7UbjBCIZ/YoZ361gpIy1b3Be2OitRnjTKhuqSfEi4ThJKxIs/mXHIK
0//5kv99ClUvoXcJinZtP7vVdeyXfzezggKCZe4swR+NDCHpz7mYEM71iqsmffltKeHZaDJKLT1v
ICjmNCYsZAI99puQ16VuN1W+YrYVR0rrU3hHkUmaG6ogBaS7k4gif77l5vO3IZzAOsOVVqIJNTo3
hRWeIZUhtYLH69CNuqewkIMW9HfhKHRI6PgjHEzvg4xRKyt8NlzA87lD7QRc/kFmQ3mdPthl3Uv6
wCaEPinm57AEa0WuwReP6fgZIJRhEXvnRwZxkrjgkuyEVXA/B0w9qhiqvl9g47CcoeYMuzq6qZ4z
ntvr5/At2QZ0VQBAHsKp3VoFBDflGv4OvwtxEjx/vCMzJ7a1N9BJGuL473eKS3SNIgrugM90hkYN
2O8Z42sRaANnAic3vkHeDsEOiTsaAR1IwWapj9HQ28D8IGfkwRp9gH90QSlvy+gWqW5L1G5aDZt+
EIneSPz7u+bTiQ2XPj1s18OCVpeEG8aJNzrFdCX1lv2gLQuZz8/CmFqpXbukB0k14itcqhjrnKjd
lx+aZ/ic0BoNAlnInBG5V/kfwmsuK5XHk1EUvmC6VsW4N+IzG2N7EyxyJpDnYzwlGU4qJ5u9BM5V
kCRly+WeW+Jo6OI+6qwmAd+GOvYdYeSA8tT9rLbqyHkUbDXIN9bExwnYynAQJZw2yoDkNCheOmyu
558B1LR4P2l3sBO3DZ+b2JAPyB+jRZifOKCg8Xmf+YgZsBW7wWMu32QwIMyfJxHhfOv+5PIqcIn0
zTeWvC+JQzPY9kOInlajeTpi7XqO1GZxN0EDcpcNlocGBOO7EqBWlAAm+b12KBYzEi2qyz5xCeSj
TPtPWFrMM0ygU8xucQ7MoUg67t1umHSHBBTUG2LULNFyeV/zPiU/siS6L+BwEscu6H8DuPdz/GiZ
KCt/ZjgTmKpudzF2wDlhER29i3ltaZaG7YcRBFUSYDcucJFQqmBW5oJ3+xTwK8BtG9WxotV4IaH+
4tiki4e674cytVFsV0Scbz1AqgH2zU1Y6t+2FTjjmLNkwT+iRZ3cq3Vcr3kSPNDIMiBYXjBbKqLY
pN3rBydDhOz6i2KSnENpDxdQcfatRQXRQ5ROrVdomxv/Y6URBYFIFAa/fU6F7pDIeKChG163cSnW
o68M39aYVsdmsCaNSo99Jno3u9F+1GSADR0dV0iTubRHgwJG2w32VGOBKcxdHVtCkLs6y1z5Wnpa
zRGtUQk2ntZUr2Rvrf8Cvqd57l+4Q+y+4VqbyeCgpRnU5+PiOO6VfHHUfqAVnMggFy3atup8fF39
orhHM6QdXPCzafsboYWsU7nI4GNfdWkwI3asL46ajaU2XIYC57PBx3wrUtyrJG5/MAt1Z4oV4K+d
9X/4I/nd0w5RcUZWdBfTRj8CS1xfA0EYYBI2LzX2hY9T5ZC7j3eUs8peO79o4NsFbWycd60uJre+
IlH1VIeNaropjbcwgY/zQri0NGPqfjzf2tXawv+U2sTDXUJooCgWOsAdLUAvUgsckmXh0a+VmaPa
RJrX91kcczGY9uHXy5kk2T90JhZmqpwgrHnkqDVKWd0qu3ZXJD/cCeZLY1V+33Wg6cDjRA6DIoH3
ik1SghKHUQ6yBe3HzUgvOPJB5udEfosiGJSPhNX9kHnFnX6CrQxOarq/8eW/W6RW+n22GUvkztgN
wArekwLC/2wyWX7UjiPHRICk4BFsfaL1H13wa8YgKgqCbeYeVAdAQjVU4JfNMG5xjpOm7yfAtvaP
M8+691a31pC5kV9fhT6giyzMJrZg+5ui8gco1jh6Gn99J+UcF9o9y2THGH75pjnuAIFhz8gcOgRD
EQLe+cWwkBFNXwm4oE8Z6wx0oZVTBptHL+QxyyIXW0okj8QVxY0Y81kTEKtrcdHkyHKJ4Xrf/t/z
smuaLJRWVmVmvR7rugg3kEJvAoSn0W4S0+3N1K4QMj8Yf6DOgnGmy+87NFF0Xb2TyLIPwVqsyyaB
zIlOZE9ZAuJexYuIo8mQHd3eNmrXQIdVqdy0F/0m88aedmWjEUhAQ5kpLYEFAywzcP0x5g95+bbF
gnyEFkiKsFRr5r5gU8AEOkgXFwZ1mCqoq0beaqWRZmqYzzTCxkHkN2B3hCkVZNxnhkfqg9DrNuEo
hcNFvh7GrJRm+JZZYpGT+rGwpyTwbbmoPmCsYZ0TNumS8JpmuQmCmgGSsaJD0HxH4sbfB+r3lIwS
DEufmUXAQ/p/HxIF7s/ob/taJxexsWODMo2f049/x/5RTWmYl5GUGKxa+SrHQQ1GF73Uvd/sfR8u
h0jd/3nvUBSgZEwd9VJEbVwf6NzfOl/UtgMXT9AK+evSE1682Os29VK210tiR3Wtp9aCcShHdaMh
YLspcL4YeYlwPjTb0vPqYvGgcHZXltfv0Jd9dVVO6/Do9MURQ3+I/no9ALhoy5kLUAmRd9fmMOdN
IU+9WLev031SfCgUvE7oX5NaDOrT8OlAQhPO6ohtG3TtERJBk83hmSkZHE1QI4pkB/cUh9ku4QWL
jD/0QitxX6Vnrr82phXWJsFMfJvbeFcmkCUNXGGLQHasE+UFgswv6Z4Gg6kJZ+F79RR3FaTVa0Ei
5rBbIVvFsamfXD6BFGkpy+ZRElSRhLjhug79KOVnyt87mEaRF4IkqEnBNme/lXRJJkb7PMkdg8pH
0cf+yPOjGH/fKd39mmaF3sIVBY5+SmplRF8C0xLyfltK/aimxaQx93BOK+iiyne9S7KAKk0yss7n
fNcv2xdk6Y8hJ5apfK8GG1iHZ5iaJp4PHbgyiNxlWO34yvhOLj92qbjoDPV0PtIo/MHdIZD5VHi0
wwQOtT07v2RmqGyNJuCJWo8KfY16Lw5tWlkDKjVPZ4/31EZd9ZaIXMRGrkjxJYOVqTdIKWgAg5NT
9NivrIFoYszl2NW0KMPg4Y9NaUcABP1ExcbMyJqbLXj9lQH6WXJfMjqZ/4giPYWyCN6QvfwFvFOk
bsp1yMczY3N8to7t2Wc+RKiTFXYi70HTLYTJO7jJ0VgW/5gdea5WovzDGzJgzpz7p5ZKKRohggYR
UIxxS1SCtP3tkN5W2QzA+uHafRBZer5ofACaJ2vSEcnxHxjlDD3Ch4P3okFAjOcfIqYLDQNZ2eHU
YaB9Q6zQYaDf8yaULH6gBB5STZMB7b4GncH8fB9+qzAc2MGSPEn+bKlB6vvNovNhxTHCKwZU4teL
etyN2lozZI0b7hTFr1NbahYSJNdh3utkAvQJTcTMPTtl3t1LcHUyTOtWJZ6uwlu7E3zbvrtUb7EK
etrGJof7rjlD4c4XP99IgbjZdNZ0eEn3Ge64URMk7NPeR/9BOCmqgapSAVm7DHxwrNc6Wp4v4qAl
7KFVK0mxYUv5qTPe2hJPOKKMjbJH5qLm4z6mxvg7dSyA1i2tz4EdNKeFSPnyedPwGnY7J7DDtZFR
N6nVEe/xhfZE1hUmA1vFFVvcqN+jX6BHf0HnTvvRKMA5RRqCjpdmDKwjsruWndyXQaSkCKTgzW8f
zrv2N2j/oV7PhZf3v2mOD6amEvig9iIvS7mDxZcmQ/pe/Hi7Q1ONgAhiZClVU8loJ8gdIjqtOiGO
jdx8g4h2JD0YjvjvAeYKT7QPvd95TPY1HJk0Mki280GVPMApW84oe0tHPBFModi/lVA+7AFUnjZL
ZGdnNrTXn1qSE9RAV+P7Gg8Obq46ifAVneeHM8MGIX0vMdcTJnSnUS6w6hjz/lQb+TK0/d/BQ135
0dcWqznm1es7oTKGxPZEjTYFr0wdJtjdN49Fd9Us0leoBaCnHINx8rhqjiX2BuPMLzzGOXNHdD1Q
UW6/YDnFpFQYE+Ca/2poS/75NSwUAJcT7jTi3sivFMte36DdHtTNcDlDvYdKz7XR4DtFmXgeCCUA
kvANoEUWFMQ0UkbfN7gCcJVOfnRANgqLqJjExDiSUqnjAxMpoQbl24zq+Pvk8C7Zxw0mzpEhKfXE
K5QsBFRjg2e832is0HAmeD4SHhZtpK8nU3rherZ82yelOPZTQFh0WhZpPDtXT2FUiWG0B7rnP7OE
vw2UVdDg0YeL2e/gDiUG7EVD0GKncToWsoY3SoW49n8FlVeBAtuY8z3M2WJE59WNGli2mmwCd3wM
G1THpPyVLchg+XCwP2D7Rtdozm+xec4lVBrXQAPknrJx/KxcKLSGLjmnYis9Dt0/mjNc8m8/uwt0
j1QW78kRF6gczRDd0hJM1zSJ7+NUH3Z13T8rWAkJ76tMOygP6GLe2eaAgSCXlYM5OZJ74W+5fTfG
sup3l125EFNlAwxya9Q6VNQzxu02y0i5D8ux392gSuPxV+Fea+Slhvne+b/pfFhINgywI5/xJZsp
+0Ar8dU6Wee8xlXToj8NGhEtiUYfmLYNCQvXFdB1fMUEmX1bzbeOLVccUdYljQwNv7ju4otKJGcz
c06YtUll2F2JfmeeglupbMYGdOv6Uwdr17InVu4UUhctzIMID5rdi02NwCXGeQPAHgiaJO6TFOMv
5V2AeB9LdQDKzwS8OxD/VZcejgb3GBawtErPSg1L3rMOUy5E6g3zN28SryPAhL/FDdqs2/ldSt/0
4ezX9RucLMLto+uoMq0F1f93jbkQpTaycHOLnl4NR6MvOjzVkehrWR9KMqNFDYqZE0LPkMQ1ww2E
JR8UQXTqHHte0f/XW3J8aDol5xRfc+5OqfFnFGeNlyCMuatFh3OvfKP+MNUcHt07bEMqh/DD5mlp
ioY0CrWfK/N1t7NM2xw4qQ8cTa0aN1HRqRfrw7Cw8nQ9FM5q3djoIlJ9fQ47mAFA5G23RiL+dima
MwstygTUKca28Mug0WLn99cmuUDBS1QgoIcDJHzESUcNqtup4Q/y0ZuTnD+08V2HWqLlfaRUtVCl
w1eO1Kh2ZPkHr9Yst8RGWoPqrUYVGu/7FHMNN2TBciN7XymGWQ/D8r5uPXiF9yaYIyYHwvs2GCmF
IeqkDClRa5rnQRbLMTQXdXc6Ps4yyxZ/XvgM/HtF1RyEJ+OChtZ4RE8d0H/UkKzHKebXLM3sWulh
38KaTV1c+jhNcEWYfyTgUN+rCx2Rm4xCdizS3IyLFMX5QvveQ+UZWwtPf2plGx3oRjJaOvsooJhT
X4rGDDNIhUu2QVxjM+PQ1HsAA7Lo6Bq/X5HsOytIWjKiM7A2G60G2ASo0OpQDMhaDE6Ab1bK0fdB
lE8sQBidyFCweaXK7qtufce6PvxVufKeKNglQxeMiePaSWnOCVUPCrj4AT3/VQscfkKKsJDj1xo8
LqhZPpO7+IOSMRuSceoOvqZ0Vuf9Kh75A9x8pHcz7X4u+8Y/+/hdJquy7iypM6ddo9tDwKOsxzix
GzBmP3VRfOGl6xmTwyB7G5jxDycsMNudm/103ZbwF3d8a6nzM1y8mmfaQ8JvVgLyY4ri3yqbkA9c
Gj2fa822SGch97bzQD1VDUnBskc6bm2Z5jf4DYIdcgAgU6odT9EZnxRC5u4dtvQw5hUa+ABsYv3f
SAR7zOrBPys66JCU+iCZmkM7LlXMnLsQUZ6EHQOSrl7g7qwjferOmGeRW71ge5W0BB/guTy2kFbj
4rkE/9RygJClTzjg/1BVKkZv0Jetk8ECwlw5eBYDn5f8YYhVfaO8REpBi/zp+LP4mTA4m1lsRYaT
yKMgO/xIN/tLOebj5muDb8khTEiLuJJI3pcUYKnKLUoCEBs0mh0cS8pgm2CHawTHDl92sqPEj9nd
Tf9rU3ac2YkmZnHJXBH/TkoS1Enr9DY3wRdUKj28Cy7NqcG65HcdeZ+L6Mo90nhZBbsT63P/E/jT
g5XZWY1OaAo6Xe5pnYwlcivTRmt9DzmCDeGzpcO0m6DoOQc9hjPDdWm3Op8gEl8HbNOKTKKJKpsy
9fpUnuzpDnAU755goUmK2mPt20DnepzaGD6MreD+lIN/cIVk/l+0BCAX3LMQ9/U6KIPzuAGBN1L/
l3NoI9AXwAMXq1JIZ58TOij4rSHwGd+La5sVwzpf0bLRptu8kIEhV2jthGijiv3qd0ndGYoUroL7
qWYDgiJhi/OihsywSWNytb2Y7DccL9bc2MqiX8VABGxAqEmHUY8yHxwEPBYxoHEc6EHBn/Z2jryN
Lp/5adNogr54I75zQGFs2Kj9gMg/jUSkt14ksSvzeLwQtKtOQS3gHh6WJogOFgrWMLZ29lloYw/f
y0yYqQ/K5MY2wNB8Q/efSLg8vhzOwfNDMfsdHHNRa7QOAjvC+oNFhH5+V6iCBmJERe3KtkQ6V3sN
nCIt0AO91VBZp0Q4xwpCBzwO2dWduNStGaBFOupCdPMkGf8wLe3KTxqBDwgvutzesCvHby0Vv0qg
RU/a1FEnm8ZjVLCNLZXQNBZjSUvPMWxVEZ48XebixJOdxKrLttM2Byq4awMLlIqC4gXsb/2sbUnx
UWdA3xbqteYCPD9Tk6eQqqR0A2Nyaz7YYTfxA9hb471cwmn7ZmeX7RQUA67QWvV5wIbnHPZ8KgY3
OeVphHaPzuvE6txKArKIN0Ch9K6kN2ncBobD7G7ZGASA3ngC61P2HXuAo04agG/62QnCheHaHypA
0CW3zU3aQSgdA0R6+0Lj41+7x3kjCDSUV+V+T1zplN+s94HoZpo4AFl9W+ecI7Ewz2uwGK/QUwQJ
ZvEFN4IAX2rUOU51IA/bxeA99pxGsQ1XIK7Njj52AGo+3aQhmqX544O/bxmPjhNwmswsf37PK9Br
F2FWsAGb91oSEclOc7loyvSK2XO9Pgr35aR1tHvCSGG/tL90f7kX590sqhSf00YevfbL0L6HSDd1
tJ+Pi02nI+56NybKeRzSZY9dU0TlkmKxh09JH93O9KbxLp0tpf29GjRukUykxhJYi6lDaxKGvoP3
/IqUN98s6kGthjqUp2xTp6x1Hv7IJLDBhJJ7bD6NRY1nW50lXWGzeBRGzVzXQ4Q4oub7MZBOr+2D
9UNic6as7zf/w79xOmQMPKhEu15edX1L1MbyDmq//PEEQl/7cNKxPNmAL4jPxxNBJzyJVFAn+sc8
G4hUFvARXgspwEeQa4RKWUMRu2L2IbIJgEyU3sr/QmqwWNekp8b8KKznQkUEL1L5q62wc0FpMLkr
yBHFvQqYTr4wm937t4PkbWalR1rjlr5IwaHK2O4sq+Yt6NgrKRf3VKCmNzXR1GVMRhE3umsJMq1S
zXAQ7DcXWzxMFwWMZGf2A7qHg8dhwg6RLqYL7ADdUWePqcSdjJChoOBor4puV+nqMy6CDufuShCw
pUdgtBw4e/In2j1or7NmoYm2iEGUbnpOV6P/Vv7YqqkR4t3nDa9dm1Hd+ZP73f6akcLSXa24vgXO
hBT7KPZ+zr4fFDoMQSebnS1UvGg+a+K8UjHr4T5Bck2XJEgsBbX87IP4uSBvzwhqeOW7pWA4WMIq
yHuxmxJNwaRh+Mjy9ewG5GjPzhVJlboKajisZG7Wr1MgfORc3pO0rLoxye8kpCNlvP1zv+sE1MuF
+9+SOvl+f1T5d0j33D5+fSRHdv7juQpY9dHSF2DJdnAC6TV5E5B5QkDh4d2DRlrlcN4EjHs9Eaig
H6+CBP0qdDZTf2O4+DITfVOj8oHjDMnqijHcYAvx6z1zZQ9fDAF09B7Z7LrOtBtAgIpFUGPxW1ZJ
TCPlswWQj+51if2/0V3umN/ppgq7l0HdzpgY17CkM46ofhrgiQy4u9eUL0L2YPsKg+Y/9O6fBYjR
+BOcUTpDGmbhG/N5IkKe5AphEot1h7lKTwnbJEKvtOcR5s8q9Q/hl9IW8Mqp/mKzbgJIu/HDLJ9Q
YRI38GISTbv7vvr3YNnLdlpeJ5owQoKmbR++zeLySSc6vcixpLMi0gYcyVCJW6zweY0LiFs+q09Z
vvuyA0YYDyGToTQhQbdwFjAXOxIyAP2ZRe/KQ7iTbHe2rK2ApgJN6nD/QdYTUvdGW3tqR4fmIE0I
1EknVmnwMPkkfWSuF4izMEhrq7kmhtshtBvg4Ro9YwhesZ+M5dJZgC0PJZR1QGb/wrCnTjszpPlY
1/YdgOqKSwCeCOFyUeNwR1q/83/lwKkh+CY=
`protect end_protected
