// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
aFmGA7ZYA2Hh7ksQ9XT09DUrt5XCGjfHva/+OhnCGKpHv1QZWWjcNiVFGp+EXKVPFxPQ7tzYuHdd
/2m3FN40SPwudgPqb9iVdfTMFAFyifrui9zvV03nkJZcI8qN7yAM5bm/lurKzo0foyfNi7+swEm9
tD9q4Af7vKc2+FXcUdSQ/o0dbGy11G5ClC8uokCjg7P2PTjLMBRjGFa/n5lfCI/m9fZXKND/sff2
fmlM+7yFvyNfTbUmlVsYWEKZl6RbvqYBikSjx+83C/xkrThIfk7ZpzUzoMnCUYBUzGHvmzdn8VOb
TIORQpuRlbSa1ZPgC6U91msPiS05pDVne17ekw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2000)
VihYqe745STTqyk9CM3OfrOHJD59/HLYRF9SWkrDTsVV0guuHb9nKXIw+N7H5KWjNesE5CqqBtEU
gg9lhd1FF9NrsUX3zpjTfwzz9MTYrG49+qIaQ0mD+eRSSK0gwfBqwHaAkCKHrj02Njb1VgYNqUSq
MUdxcTzthV9N+AYMveQDWk5hzfE8VgDlUHEvUpCZA69kYddhYXZvvcfl51h9XJZFfCNshuF9cmMR
PK92K/uPnvAdAkGE+CcQDdQ4Q+1rIYgT4pyQaxrNdamf9S709yDqV16rtJVEQX+PmTcWCcPLL+Mc
0l7PF01WoNboA1z3CGTDLXaNQntQlPxooNAZlRM5ZFThe30s+hxwv/lKZpAbYuqk1Dbxzn8Nray+
GhohCwiqJ9f+Q53uOB1AN7993sIBSym4gpiS64GUrAZIEG91mN7F5dmYDQipLBDFoHKAUQTvtF67
MCCZl20LJE0fwRBSlVESJFbzVviQtnuS1pHI2Q0Oxp/LmgOrLsz3tDaAUYDi57VhbIJyXckAEkun
kuRoJrIj2W+l3gQWxCbfQLMXtxFY6awYN59SI6rG/lxk80maS8pONzDuNRFQCHgKDmaFrloh5Cj6
qUF9llq5RZp1t3FcjuihRHqdeaFJxaZFInUHv91T2ITHjoVe2blKysa41deCDteb3W9GfLzwWu/n
8rP7FM6QX9qvaRE1w6xUG5G98F3AFhfGpZqiXqKSC3pwCEJ2HYmsvnF+DY4frBxvwQMsUQkfFi72
8RbGpO+A7wu1encQjYlYutd9GOWFAWcBtUCpfuFlr6UUvqohsNeoZ5cF312IZJThuJQRfVJQpfR3
72sliaMkW1T59Hkym1mBTEa5bHf0letH0Ypt2aWeuVtkM/lIlYVoacwwDUN3G/WQt7S2lN5tMUSu
FZ18LgYYCaqoUAnjXshQIc88+Kx1KhZo+zyFdOuQUgf7+xf32lfPRnxPi7WtWAaygR2JRMUvu/x0
+JFsIcW3WEz03EW77AcPQodOkB9Bv63TR629yctD8lhg0IVQPHRxGB5imAkODTlyVnoo5EoWADKD
qaCb3/bqnPa1e/1A6MF2QQ+52X8VEFVedNdGkb7Ggjj4spVduMAB0z0VT+CoQO9DvB/Ye/5Ji6to
+IDdkSdBLLIurogl6HyFIQSBCMtWGgSiBcNacPXC0b81vnCDO8yvWN1QTBeTtM0a3wt2MBa4Qpnf
qjjoTteV/s3jEMws1VBCplbChBEp+goPDm+jM+wGLksSy2pgstSqwjiEo+KnTf9Mxi5nr2j9+6Ef
Ja9Ni6eHJKxE76MWLHnLHLaYTylMOnn/5TnGUm7spNetwVhue1rKLLu6G4MlqZRN5yyiGi+lXPkc
YrWYdG3z1dbqxkyfzCecnvMuClLSvq8y1vJOPN1ytmF4qIm/3YJwFy72xTAULkvO7fc8vr2Yfncv
zKgc/yFWW8a/0X7yVmlnLCCUtyxSsWfJime2OmtMIuX3AmUpszztFuLGg9JWiausK4V3Hf8H7O1a
rfb65emuf/+rIdZf4c0bYaV2XLWV6qsVbGYJc01lo7PABOQydgL0l1wc8G0je/zOZF1eDtWZ1Pdm
w5tyxXEr/97QDc6JzHG/h2OMfbMLl4+EDhP1QuaZyzA1dkTBpY0xYF/RrbDS2L4c/gBHpaGn1swr
Ao9gyKaE9Fb2XYCtFeDGx436DGJvBOhg8bWw/XIt054aQS0FHDo5xX5tAXdaocfcEGPe6PLCsszJ
yFK2I7TEQJINWZwLIRpv3mYq4tT7qpkeJ5Z1aogE9idRYDd9/WzWsYnVffk6TV3oIO6foqTpr1MG
jsz4HxHZi/dB1LMl2dKbRL/kYHmduDJQIGuG9BrHAncIPrtVNZWRG+WMO+wZp07g5bgmFBhEWtK6
iWCGWWCGE/ycfFJcrWkeSrPVI+UdFCGgEu2C55RC5wL52b/lktkFHrr4nVpYBJ0/Fd1JSJ9fx6cx
zHgCib3zhyn4/mjkANS/Tc785kikou0v2/uE9jb+NxKJEna+LqXpgPyu6a0qDh34SEIahFY4W9Yn
uQXZ7JUgHrAEZfgBX64Gv/6fNHCQn45ldiUn3Ka2mimj637w6YAuCPRn4hbRchpGe/YhKg87H6A6
YPJdSFaTQVItwB2qImKgUFyWzvrMLwyQMrcpCL22A/MO+WC99VPn0fgyuIQZKFQonZQGCPvG4VtM
B79+XNnZ1n0BpbQuaOiqPLbNEEYIlddz6fQVAZtmrSeUms227jpeQwrCk2+1/MUu0YM1xRhjTmy8
TvVdtj18bDCIgqlrcLsL12GpOL/jIf5h8mxHXoSGy8lhWSmLA9gw1koBk/5c9aj+fdtXbu4YFjDC
Djgaf5XtJBTN0tineJtqwADH1wV3nkGA3hDEn2IrlOfJ2mm7zsyr8z8S3Uxem5OF8LjlIfa48dMW
hg1SO2BEAO3aZG6HBWMr2KvoqcUy6s4h08MrVbt7Qh+fFQb9JpQTLYFUye81w1+6eyX0HDgobn8E
my2Oo2logZbSv4S7f3j7JV4T5NVPMWhMJ5kjU5HVa0ZBUfmyQV/UrQFevo7yYQBU12IgH/YFURTV
2nx6IT/th9OTF0XnLjjArYwiy/xKd93kieYxCxtaoYR4ZNj21P9+xmDd/vsJ4P37UzamPNoqsgdW
IcOhzDQ=
`pragma protect end_protected
