��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[/������ۆ���
�yB��UR�� Eb���ub�j��V�
T)���	K�iQb��F9K��[KOh����vr�� ��N��F�n���+ ��H���{�C�V��a��p�E �q�>�(9-(��_��NXu�E�芿٢���n��އ�.��T����/�lL<;B���AwfA4N��H��b�6�"飭3j�I^
��H�M}�ѣ>�]+�JA$�ڻu�G�Ѣ;�u~K����z�������A�QbC��0D���;���s� ��v�Ef�AZ)4�t!�ug�"Ku�Xó��Q�%[���^�dyӘ������[��#�d�� ��	�\u����'oi�g�V8_G޺/�U}��'y⵳�P��4�_^2���	B*G�hn<�a������K��������-Y��
K��®�ᗾ^�n�S�q}Y<!��R�lk��'n�IW�(����*G�~Wm�[����iPn>��>g!�C�Mه&>��'�r�M��xg8ٌ;�r�@Oy�[�ò�@t�dB�b:���=(�}0�2�T?��­��뻍����9m5����$͌o@F�$�6��t��̓֬bA]l�3S���G(�K���H�kD8��d��hF�'�j7�c㽇���)fj�X3���7I;����s���&��J$�_�Y�/ǒ7��9�Ї�&!p>�7&��L�bW|�&¡M��H)8:DP�!P��ot�m��]�O�&-5^CV	�V�:PDAw[e,YjV��.3�b�3�,'�4���5���e�u�-/��G�H�,��1��p�RE��+k�q�J.���	Gխ~u3��')��׫��X:B_�Z#�¹�������ڐ|��B���-�I7;1�����M��p��r�29�e����o#�p��Lo�:�b�+gſB�ŷ��OXP!�I`=�Wv����(��Ȋ�-�n'1�9̭�<uS�d��Q��t"��R�i�V�&�4���j`�xy��/�����+y�Y��K�t`2���h����������Dl`.ҿ��݂H7"��]�WJ�W����:�oT8{ʈa�L7[ŧ�;2�XD�
X�<�L�nV��ήF�f��.L�RN��s�e�q�rw�f	A�����A�(PV긆�;�a�ʐe
��#+�l��j������~�2k�Z�Y�ݢ颱�d+�ks�rc���1^~y��$*d�k�0kQ5 ��핖�\q���X���㋍�� DP;^�T�������Oka��"j��@��E_��8|��qmu�h��{*��JSds=��.!������9q���W��á��	��*t'�}MA���֎]����A$��C�W_;���@�xA͵<.�EP�wpv烑J"JV��'���@���U���^`G��sФ�R���?ϙ����Wl��~}���.�l��3Q�-+�fW�����)�QT����J�E�Д`�l��$�ڼH(�z�V�Jz������H��<^��e#�o�׺�1mo�b.�!#k�8�+C\�'��L�I�;�Z_}��(�f_bu`�ff?7yCآ�àFS+�)��w&�H�.����s�/�k���5��T��L%��lhB�ҵM���d5�io6�6�q>�r�G�!�ީ�2�F��6L���8k��3w�"	���ND1�]Zn0����C:���'E�w�s�چf��R��(�!85�>S��D��?�y_�o��y���RP}����0Q��BUlŪ�bO��=�c��}$���ЛAF�a~�c�L�oT��G����D�D��'����F�l�O�!l�b���I��v��	�L�
z�YB�b�ݮz~^#���sو�~ѵ�d�7��>L�ϧ�{!�AqW,b�}��&2�	���'�,��skh�ׄ:��0+��g�Pk�y�A���{��i��|�e/�cMo�5�h{��m������* ���:i6����ƓV6����sǜ��іfP2��H ��i����舽�t3n�H� J�.���==H�-��Zt�*�F%��BP]���`�%��z)�.tǇy��X�Qq�Q<�R�z?��8 �uR�j=[W����S�uZR �6;n���¶<!bd��$�tH�є�qK���`��ꉋ�pW�C_�ь�)H���3Bu·������c��z��+"3*Xo�;�Q"U*,<�}����V��g�����������8�|?�q�l���
$GH㦸�ʹ?�^u!�����9u4 {��F �����!�8*�D���Y|���^$�ڤPI{�(���n���L^���T�e��|�:����lq�k;���=Ԩ�+P�;t��]$�IO%a;�'7n��~�u'+�P��u����¹�lr�G���p�!�$�?Y�|��Z�vޞ�Z��59��~�l��L��<�K��C�"X��SiR�E8(J#N�_�"+h� �VpY0���ӥᕴY��z�K��u�N�J2�����tEӦ	�қw��2xiJc-�La�
J�N�׶>+�[ ߯ғT�S�z,兙�au`�-�!����n���J6�W[Gg���4R����U��.7�\!�`��Jf��e��m��Q��7J��ki�oa�bQ�1�������C��`�KU��A���"�Lv�a�vB�|6��sP{���.7K�/��o�F��Ԃ����w��
�:dr%$�(;SA.)��B-O��cM��'�H�-����%��x� �z,e�D.�m�H��k���$S�q|o�t�!��Y�\Yv<X��	j�r������R�Eg��!{t%�_����h@��`�#�Ǡ�Du��VU�9�c(a�3�`�C	5�I�2N��8';�x�4.�����e��ɟh�B<�n1F]>�65xg!�"O��M��iw UĻ����$��؀&$��QP�a�I�c��o�V3c,1W:����dbE:��u>�����p�صd~�&�1�Z$="��-�!��`G�#��\u��ad8Qb}�A�q����Р�z �}��K1K�p���,1c��X�v�ώ�j� q���W�N����\�L��+��l7inq�O�̈B|���o�M���0�F�Z�R'�4#o������ND0����66�t�,X� �z��q2+[��{�=�YME}+ a��Y_{q��<�O�B�C���V;�CI���h�Ia F �����j��=TWj�B�ui��/�G&3����oP��qP��G��G�i�|Q��Ҥs�:n�x+�ĩ���M��c�լ�b`��9����o�Q_����k%�V�3{�b��O�;%�nj��Q��o��Y����ϝ�Եm�t$�ٛ96|RM7j/�2}fD�)�'w�";K�l>Ւb4k;�oH��0i���H��-T]�Y�M��CUaEWNMk�rĚ���H�;�����ь����e��v*s���jp\����^6nGL��(P�}N�+��m�����f� )g.�
U
�>a���X����gr��x)q�H�X���\��%��oz�H��n�rC�PK�s�a�$�݆�J�S�(ptr"{Ua�4Ϝ�C�H���q��!�z (n��0G����0��I������m��'�|�PA�0�X4e8�e�"�Z#��FB+�Q����9���U���9�1�8 z��V�J��~�]7ӝ�ƀ���S`��*9wޚ�cY_ g�u��ebt�t� � �s>-m�1N{?��I�f<ZݛC�_�W��q�*�B�������Ѣ��xD6y�a��Y ڃޏ3k}@�Ҧ��*��������q��y|r|_p)+%���FK��)�,-����̙fu����!	#@�F��xq�7�;�L[��=�hc�� ��Oy��l�����B��}�Gӄ�����i{�o���{?zh�u���ݮC��"�����s�9��تr����ʺ�k���/2kM�V*��[����Z��%B�5��J��ay�FE&���s����w���b
G�V�D�"�XG���:D0��������$$[�^��e	Ƌ����/��~�1�w�pе�qs &��1�Z�mq���Y2��/��2��U�+!�����8L��>�H��cR+4lAЖ	d8:yag߼T��~�����iD��ա�<�nW���и���Ń��7f����B�ٕ;3U4-dCg�!rϸ7�z<Cg�!�0�n��&W^%Zs�D�&����"�`S���Q��!�K
ǒ��2�I��ò3R\��az��(t�W���X�:Qs~���}��*��lUu�X�x�����P�M���hL�c
���}Y��/�N]i�kS Ʀ6��t� 3��c�����
�h�>��vx�]���1�P�&��4\�S�8nj��	�u���yN܁5�� ����fs))���o�8p�8񴤢�4g߅�V=���
�*|
�ӥ�B ��z�!�_�}a��	A�S�o����_�";�G"!&%�b��bG�qB���� kJއ>�5�?��	�?�t�ew�ZS�C��p�	)�� ��v�A!1�p
>�Z�Y�-�v��*�#.��R��ܨ����QS-%.p�����I3w�6U�JTt:;�+ݤ��+�ȦFulX�o�w���
�ZB�j�$4�K�����������}U��:�#q�AR�0�y�0��T���Hr��Ϭx�if�b#�)j%CȀ��/�b��T��u?g�C,�Kǌb���5y���k�ge'9Y���)�5�>$-����k���F�g�	�M2���9��~���o���M΋IK`O�z`�RK��G��}��c�.���Z�:�z'	0rEAR+��*����E�wO���[�*���./,�)���R?���E�e��2:���:���#FҒ}��r��$�ʪ,&���y�����>��|�;�X2�����P��Z:��h�$p ��1��9��ƺn3� A%�~ \6O���	'u�B
^%u�(@��hr�����?��ٵ�9�}�����S�H̪R]Q��\��/���l5���4��G����Jhw�ߘ]�,��ڨ?�8��ƕ1gp�*ݛ�$)�?�7^��˸��(�l"QșQ ���ֵ�;�c�s��h���;M)?���%������f� K�ev:>Z���v1���k������b���?�٧;��V{���4�RXf��S�
��s�N?!�A�]DR���e���q[�'����ʴ[%roɵ�F��Yl��6�u�����C، 	I��I���͡�����߀�ÈJ�d��[�N\W/Y��F%�k&���}����@��6�/�����":	����O�<;���zq,.r�C?�4d�aTAc�r4Ҟ�����6vJ�hrߤ{�=�5�5<7V۾�#����@h�q}+x��=X��3t{�Q۟6̅����e���[�>��d��9��Y��=BU<�n��Qx-#��߹�O>�Z ����%chq%�p+M�Z/�W���>�&�7�S@�I'j�7�M/�;Xy�q	�7�ӣ=�A���{���TSF���f%���cׁ�SƉfٳ�!ki��oj|6]�@)�eL�]����.�����#��تa4����{���M�m��t�5��T�ҽ�9}J�sj�h�����|	Oq�ڻ�ŶJ�E�O{
��h�]⇣v�,�&���������l���Mb�7�D&���p���>�� �)=s�#��(�đ�z��q��^#g�O'�"*4�?�1��h�Z�5��2��.IS�Xo�rYb0h��ke�4B�>KT 2=��b�o' n �M;ݨ���A�������mx�@ay�Iг��9 ��!�x%P����ܞ���`,���N��2��+1m�,��#�$���l��P�{f5�*�q az����t��߉U��d=_�*�0�]�4؃W��oփP�n ��tơ$�����¿��q&���l�~�S�4�%��n>��-�I�A����m���$~ܺ�\T{�1����m=�و�S�AA���:�EJXW1x�ER\�J!���|�s�  ��������2���32�(�q/j��'�V+X�h߲�PM1X5��c �Tȫh&ܦ0��]��dy���#V�c�2ѣ�� �N�Ճ��%,��Wf�I��"�����_P�/ˉ{���-
Px1��w��ʋ*��$��z�(]���A�1Tŗu1���5'������P��g�IJ�@�JJ�	��iʈe*�5ۀѩ��1!��m+q	�hg�҆I���ߙ�< ~x��2��W��f�ڼ��Uv�C�g��	u]f>&�3���>�x���L�!�!��@A//�	��*n��8j�]C���/���Y:����y0d5�O��tu���-b����#�"����Y[�s�&P{�G���7&y"ѯ}DJگA���Ol���;C�*3����7v�r��v3��Y	H�<o���7�����%�����2����\bHT���V�S�MO*Z:�/O�״�bab+��r�����~0�����c�϶|ja��,4��f2�>S���Sc�δ�z ����Fn!���:�#F|���v��mME�{�Ng;��l_�"v��J�]_�ս�{"�J�iW*6�V���B^-]&Y��% &����nX�h�� ��Z:�b��C������O7c��	`r�Ϝbu��� ��yϭvMEÔ#��w�C|���?s���l��������!�z�)��������@�+��YE�/�y<( X�]���s�X�T#�����PL��D}|���8x���[�7d�����>��f��?!X�bmmk�p��͘<�&���R�@�OZx]0�x��t>�ww�����F�P��B8\X�fmL�9|Q@��P~ګ��y�_O~���l���nG7�'IJI�Ɉ�����UY�>�@�g$'�m³D���֩�XY�+gx�;���[��#��E�G���"W���R����,% �X���ͯX�y������{�9�t���x�$�]{��P�~�[�G�e���Ԁ��vʊO`hc�;�bsU?�ߡCC�z�aAy�|��\�P` ��&��^I�2�ǅ�������Rb��>Y�&�]�i�R!&��!�ќ�|�יH��`�&0���A܍�����_I5�8���`K�`��MmP�3/K-��e��xx'�KW#&Q���aIv�$�"����UM����[�<w��?��P&��%˳��H	]�Z���݉�f�)B����3��<������s�V%�� �E���q��"���x�K֞���)ַ�Ͷ�2H����"(�C0�X�f�|�n�y�ࠃ $�4H���	.��cg����x_��'�Xʃ��C���m"X�ߩ�`�jJ�b���⌸��O����������_6 O@VvV�cȴQ7r4���L����I�'Zx}�6�8cT�w�%|
��4rX���M�ׇ@![��&�_5�Kq�Cj��Vu_v(�i��_�2S�%�Qr�k�X����>���Ewȇ�w���z�:a�Aٓ�~���p��Y�Q�r�C�v������=wb6��o���'�nq��2���<�6ǋ	�!ꁻ��Qp��rX�uP���|�� @,Ӟ�� ;�Y��ɗ��O�/7�͵�7�c1=��"�~*H<0_���Z���u�/'N �=r�C�Y���ǣqI�W��1���{�K"m��V��)���e���cN^������l=9������`��I�(��znK֪� >�Zf��̰�T��Z+m��V�����={c�o�U��,n�� ��h������g8�\,����A0�"aq���{��g�f�n�UH�(8��9@����I�ə�%m�Tqs^!Q4Ag5H��<}��h�3���!���z+�v5��HcS�'�S�`?��""�\�+�N�s����پXVs�:P$�
�/&�J.���zF�h�0%��'�{Q����8����Jhl{��Ƙv�'������_�����66�M�Oii�|�c��(��-V+03
-XȮV�O����v#Li��x�dl�)Nc2�(n�i`ϝ=���r}���W<,ۡ|�u��.Oc�"j4C�K��U����&�Z�=�)�(k# 9Э�6	0D�/S�Ò�o^m	UM�����Z_���1p��˯��F"�K��=�ޝ�����U��={���l�l�'�\���7l��У\��^�Bj��y���I�B�t.W�&��\m�q"���Jx{�Q>m�b�b�f�Oˌ���皖 %�� �G���)��֮;ٖ���~y���+�;�N����d>!$���t�N����U�A�le5 Ka�"9�K��FH��X� �{�g`O~���O�*Ґ�Ʉ�ٟ��a�1LX�"h�U�F�F�K�dS��/Eu���i8���]R�}��y�*��w��rM}7)��Zj��6�|�O~�+�H��M/��(�h�����*�|�\�>�q|ä�&a���S��nL���n$EC;ٟ6y(�ѝ�F?�Ǔ��1��	'�f>�婬���#|�O�l�7�6I�{����DQ)��dm�}*}��3��8�t��/z������X�Ov�.�ƪ��\���mgM��{ɮ�)B�;a!�|��0���@1b`:�c��c�9�\�qS���*������"t�����p�����Ѩ���n������mW�C�Zd0�%�z)1A;vIsf>��;��/ׅ�N��֖�P���'h�8��[�D�ZF����i:��`�/P��A@^�TH]�I�{z噶���a ��]n���D�l�.}��'�n��QIO9PNȼ�}��h��c����[��MʕP`�]0n�|cr��=�݆�	<n����YJ�s��.ߕ��P!/*�Wٔ埕�%;�� �k̄���"����c��',��P��$*���S�|T��َi|r���uR��hј�v*���׮����bX/e�Vi�	0�oѧl���"��G`�5mG$Qт���O$�A�ZxV������*f��ז�)���-�0%4׃�Ł�vWa�>����m�-��������u�5j�/1-��']-U�:��2�)�+���Z�Ǐ!�n��YcX���?�����a�S�і����kQ��&*�R�1脚_�tk��2�Y�)��_gZAS�W�a�҅�C�"�JX;�r���������+WS�%Ogiޞ
,T����˒��o�G+*ʹ��� ��&k׮籶r�v�z�÷�,�C�q+�ڕ,7$�K�0�n�&�9��na򯓛��[�k����S)"�99,�	�z>� .���J�K?�QHd����hޠ�Uft�]�}D�nr�u��nL�@��c#��B`�W��ʬ��G�)�q�$F�xEy�ѧ��ޯ��y��{O�#����K<Ӵ�D>�d��&�i*�Zky�ռ�i���Ҙ��M�%$"ϾJ�W�GLWՀ�[`q�f�#�fm�B!ovh��Zb:�m{`5�S�t���c���	�r[(·�SK�#G� "�H�IM���Z�u��'�H>2bȽW��K�l�J��/?ċP,Ǧ��H�%����ј�o�L��<12^DR5�t����
>�]�%0��8�1�u9�*�-�����Ʈ�M��s9�7nKs=�vT߅b��YCP�>S����%p�P�U���@ ����6��v��<\�2�vf����H��%C$���d�U�o��0��z��^>���]c	����7�I���%�l�GPځ�E������e*�(`�s"o>��.�*��4����kzc	����(R�u�j#&��oL�\�u`��g	p$���m]9a��}� ,R�'ǂ庵�)���������V��<?���ޗ��|�p�� 	̬�� ��t7o%����B�٣�!m�cO��
D�Dw�,�G|����]��f4��(L�C�v�Y@fDw�&�)��"5�ɳ�f�J!��8)Tg �7��!E���`L�/0u��gS4��ՆT�K_l\�P���i�O%�Jc2�z�B%�|�+�WjY�6�]����F��H����U��t�z����|�eQ&�F����s�P+���˙�y�^e����:R�d���$@��a�v��5a��]5���z�F�5V����V_��4\�x���[���\�F�H�I��+��upD�㕤H��6��Oa>���;N-#�=WHZ��3v�w�b�Kૐ�揲�ݣ���P)��yh=!��@1�~��u�����FLL�1c�lR��vC��SY�M�P��wn�� �#z�������^G�>T��QۋH9�|쨪�ĕq*_�Ɗ��(���v�ޚD<���z��"9t"�&6�>6�=	�  3+Q�S�(Q��dD��rA���C"|�1fF�X�(M+z�d}��詶�
�T�^~-��yq�NWl��<u��}�&:��:��ji� {�0Np��|�f��]��5m�4hZ���m0��6���v�=�2M���6�@��@���v��B�3�e���&b{P8��5��=V�S��?0�}���m���K���:�A��]'B		
�o��� x�pͩ:����ٶ3�x��q�06���BPk=�å�	߲t(��rz��������0�&�{5H�dÃ�ؚw	hM`��A��%����j@������GLek��,@������� ?��3P���n4�m<��p4�đ�M�4��<�.S��|��Lp� �Gױ)9�Q�zX("N�m"+�1F�wL�i�w|�������*����?q�i�Q�su�Y0�!�����>�s�C���1o7Ǎp\f�L��+�V�
3�P�]S��C	��gN�6NP~q[)������T+����E��qg�#���s�"��:�.�\)�AkB���g�{z^{����eQ�!���\�4�?2�!���щ�7�I�]R��d�����B,�D���@�98_���.C8-�M�O��,���.`Q/r�c��peZd��h�[
�G�T,� ���Xw[h�8��@<2�i�m�Ao�W�_�6V��$Z(��~=�P�7����`|�M���J�v���s�6���g��d�,�B���|H���W��#MC�5�lP�z�&���ߤ��	A~oc�	#�(�Rʟa�|���Ř%�J�Q;�Ӝ��}�P5�;f�c7���[����w�g�� M��40ʫ~�._N���y��,�5*��-�c�b嗍x�}�ާ�
wPL�57�s��M�N�M���J�n�r��z~5��D���Z�E�j��� Bj��0 Z��;b�#����{>�z0[�X�Q�1?D5��똿�o�ivề�B��U�ن�>匷�E��mrz�,�/N��08�{���Dԕ�ڽ�5eA)*5�ŵ��j�H>~�N��ԛH,9i.K�a�P�����f'Q8��O�E�x�Bj��K�gps3'��$�~��ţ�T���$�����u�t��i���R�s�Y��0�%$p�(}a�[O#����ݲl�ǅiR���wԞ�=fv����Q���85��*k����N�r�cv���zt
����2�3�������+TS�3�@���Ki��X�aS����v�[���Jx�ܶ���`���������d��<���.!�U�q?f$���N��nR�gς�w�^�ʼ��Ow2	��j6�w�پmĒ-~�����׈�cA��G��i��m��cA��߱a�r�n�a��ԣu�������Y�cȍ?��?-:ZQѷ9���d���F�Ӭ���nJ����in<{9�Za���af��]&��B�Ȍ�"Y7�/���>�!�.~�^]�.�8�R��P�Oi��H��n��S��c _p��ÙKY�O��������?�BW%�+lr2@�>�"Βv��8�ϣ%��#О�����P����@��G�L���8� q�駺�&�jRaQ��9�m�>pnBA�g�����h�S7�{�`�Ɯ�0R��X��B��yv��ŭ�j�Q�ν����^eO���wV}=�,z�%�9)_}�Yk�.{�4W4�8�6�(�ϒ��9�H>:�u~�.J�d������}�Vkx�[ς���#%���Õ6"k|�>	J�F���J]�mQ�^�t~���M)�9��N�Djߕ�3$����x-����>!T�}IC��[=`�׻R0��W��(@�r�~���!��D���!��=j��il�����	z���(��C�6G��G"�Ə�~~�����NDWJ��&�^ɰ3zv��+�k�
��4p�vjPRU�>���X>Y��� ��\���T��i{��7ؔ/�ԅ�m��3v׼��P���l5 �m#�̴���g�(��$ɠ�8�]�u�`Z*�敩���iV���[��:�b�j�t��O�]G�YPh����������"Ʈ�0��'mR�c� �[M���-p*0m��#�4��ʪQ�fZKlAvh�������O��K���:h��3�z9�Z