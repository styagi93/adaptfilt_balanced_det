��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[/�����������'����UZ�������(�ۜ�6yю�%M�P�������=�ZD�ݵd�Nx_Ok΅�%C�� 腤Y��h�c��W��B��l��;�/a{S� ��\�T��bX�F*�~�i���z|�s�N�܎�����.�W?�{-,=\|h�sJ�4m�:��LA��պ'5�����i��B3ʁ�I��S�S��2o��5�U�4�ܘ�8yYU����D;�Tf��0`��x,<��s�����;��V n/S-���7Y�h<^$j�F���w���f�akS�5� %\�/ё�����x���A
�f��,P'��~���rI��} ����IR��5���=�1�\'޽���:2sC�8�&A	Qm�|{�ȶmq�\i)E��(w4�H��DZFw��ռ �G~I�R7K� ��"? ]������� fC��W.r#�����y��gϸ�gS��S�0���|�?�(�qk5G=�Q���jr?EM��WEa9�L��.:�:����X��*�D�)�����HܡO������ 2��͔`��s
�Ì����W
�	�:���#����I_$ٽ��\�1O D4���e�簓�,�L��'$n��h��N>��+�}��,[�:�����fpk{�M�V�+([d��c�y\�h�h�8%�RlE�5�Te�e������W��hl�滂��]y"�o�X-���U �zE?D�ɹ�$� k`-�X\FCR��O����;*�+�!"	�W��e,�� 6�[��q�۪���]���7�e_���oF��LD�Gӹ݁���j+,�1�D�mc�Ng�h�F&N{)��ͺ���!Q%c�I��$I�����%W��b�G{h�r:����!U6��­�z��G�qZ}��F�&Y�#�M���������E���Ƚ�,�'�e��{ʶ�ƛe\�ɠ������9j�[ ���,��Dy1��y䷛���"Tѱ!� �]�I0��*Ej����2��o��_��Q�����J�պ �a�4�^T��h��5,C�����|�+����[�PQ��ٌk=-�4��8�}����D�	l���B�q�uX�U3��79����rTh��g�n�@a�/n�C�nO�+-^���<L=�p(Ϫ�(����3}�,�yN*f�����2�yـ�Tj��� q~u�̗�fw+�C�����]�3��Q����F���p�v�a1[h�tB��၅F��[���wc���b�uTخ`�R9I��b����^+��3��*	P��*�X��9��P�Q�Yn��)�I�N+~G�f8C<��dX��Νk`.(��8�������S�r(���C&
�#����Ih���Q#p5�m�z�ظ��D��I��(���Ƥ��O�f���P�$)�J-Nv��0��c��lv>�F�UW&����:#���4�g�s�iGJ?���;?�g*����q�7�{\ea�,��eb�������]�ΐ��#�N�$q�i�):
X�1�\Ib���>~��k�|�.�N1���
YZc��� ������mUL�O��� ڴ%M`��VS�:>ΨP�^}��hd�Q�3ky�#�-TVo(��S��ݷ{�������B��(�{��rq�m�lb9bd�J�m/�2�4�j�/17�ɵں�=b��� U�6h�g��%\y*M[>x�2q�r>�{H�U��ߚ�Mݹ�$uU����Nu2R���r�W��p�=��j���:�X�I�<-U��S=Z<لصaO��|��nW"n����۪�\������*C�Q��N�mM�V`�h��l	n�ۂ�ԡ���l@�#�)}��y�_��U��ev��Og��n�k�(����Y��nlA}'=�a�pF>%��_��,Eg>
��ȚF����P��)q0�]�o�ǂɭ{��?�ĐE=$����	|�6ED9`���苵h$�����g�=��OIr҈��s\)�o�f!������%2L�B���f'��9�3�|Q�q�ƍK��QI��Z�Xᤣ~ �/O��AwJ�%X��v�r�8W�{�4 }O�B����)�����ZЪO3�[u��**��A����JW4�i�qS �
�qf��s`�p�Ӌne��9j��JAh1�a����H�M38���f%���I�����ُ�%�u�ХI0ŭ��Ӷ6պ��>������QY�e?�sk�0{�mq��)����RW<�Vn&�zм�g|�B���.?����{BB��7�ݡ�-g|R�ʏR� >���E��D����������	�iV�"t�P��#���eʙ\�jÍ �8�+ �J :rK���x?�ˡ-9�'���u��[�#�������0TRީ߇�_� �F���]%P)B"x�Q�R�~WNcf���o�(@��,��#��t��+��nuMS�x�F��j��r�tn��{��FZ���X���9$���P'���^	:Ŋ����j>�e68���P������v�3�~�R\���d�ѿ��Q�)�hP��#qS�$�G�L:��5)��Z6�wh�-����s=2�Z&=���ˏ��~������U�C;t��s��yZ%:ex,
���g_��OTH�I�i�O�U�Ev��̖U��{<X� ����r�����s9�g��6��dˌ���R��3v��$U�OE�&tE-�v4u���%a'7�	�C�pj��L*��lW�
-�&^�L�A; �׉�) b�ί8�L�h����OM���ᬐʓVj�� �Fm	Z�u�ޮq����F�0�����Qf���H%]8�5���=~lD��K�s��H�pl�����<�za1�����\�gy���gp�uթy֝89�v-0&"9��A�L��Q;�2��B��¹5�
�u�M�u�QeI=J!,���[��,��[ӊ��g��n���ma��˖+6@��� ���X=����E�HdM������oԩ�L�Mh��+����M
��0�k6x��p�5EŬ��v�6�Kn5�R��!�����Dg���4gx?����-�ǝ���ќ�f�Y��kM%q��1�<���������<�X�٥|��>�
���;�A!t�Ᵽ�%�WX�g4E6�`ho��]t�Z"��K��^�8)��QI�[���Uo#G]g���i�L5�^�2���>���ĺ%��%4��ۡ���'^Z��y����F+��������i�N��m��k����~�,��(I�fvO����fh����e��ྟ0ylP���}�y���ϔ��UN�� �r�?~jyLeқ_6o"��Dr��\&�%ت����e���q|��k��-�V�Du���ދ��>`�y7����d� �$[�+��d_�T��a
�D9�-٦^�^<�ȡ��)-y�(�9��[�
jPy��!���J���w�LHW����EK��z�.�Q+8��^����$}9~�ѣ�/��B9U4!qtim�w+�!˿=�̬4�U^�9��6�]g=��H���-
*���v���Q������\1�%�Bֆ�\s-��V��tq ��B�P�I�с"dQt&Ν4YD}�3��7k�S��S�%��P�C#�N���c�����%��jˉ+��v�����!�cO����L���N7ş�<�����!��a� �Q:љ�Fv�c ̂�<���˫��x5*��$���ՠ�T֧<�w&�lmnG���Z�~Ŭ;ۋ{�!�r8��.�Q�4��\PY�r��8��W��=�JE%��u��fvd�W[x���d�Azr?Bժz�
���L���j*�*W�������ٹn��������+�-Zgq�q6� ��B�2��pGv=<��pȍD����8m��t��clEZ<8z����$��41�EW�Gr{{�Ki?��v4�d�nI�s�S�>�&��	Gv�iil��f��\�,���aH�l�y��ϛ�uS�Y�;:}X�s���~�v�\}B��\s-�ٕ�^�TM�c�.�������M6�^&���v K�����Nc���0\��� |5��X�^R{�֭�{L��R��T]��l~4�8��x��3WS��f�(��P����u\�m������A�5?6��@G)Ij��n����3��V������>��fvwq����ޫӍ#��P$�t/�kH(��V�y��䂖�k�
&���3��R�KDN�hE��ě�&~z`wl1c���������\�[I�b�T¢n��w��4Q۪r�D?2�x��5�ObY�#s4����1�/�7�6|<-�(ԕ���4t�ugS�GF�`Z�Q]PL�����Q�
��%5�_�������N�L��#&0���!�l*;#j8��@`o���E�d{���;�XrgH����ԷO�֞^��Z���Z��ԇW<cʄ���x�h��w1ޓ"�[Y�k�2�L���5~G���_"�F"o���궫��^�؇�\��,���=1ػ���0AS'?B�_u�`;,MK6�0���:&�4�!%�
�x5�-���u;������T�̅�I��G��S��ݏ�"}�2��+:��9��D��wM�J�w�<��ݞ+�`B�넋4�|�0�k�X�,�\ �S�]R� �}�7�R��y�k�c�ه5��q�9�%�.I[��$��Ԥ�b ��ղF����t~�OvN�����b�I Pܔ��/�&h�q�W{�@���%X�]�^�j�J�ϫ��8>Z5���������p^�o��O4hmZ��o#��Y���I�)���S.t�E���'H>�"J�������ʅ[o�A�@Qqĩ1i\w����#ֵӯ��*���t��ˏ:���]4�H�)nr_�<q�]H&�w����͗�.��$䲂�һE�H/�u`{/��Vw�e
�:�Kk�EN���l��]�j3�b���ǥ���Z�=�|��ߍ�v��˶.�*��~s
틯+����
�۽�����E �r1�n���l��!�ɯ��EDu.%��r���gƟq�=m-��Nz��Ɣq�����7�+���yf�p{�����Ҥ���Շ�5��WF�K�����/����M@4y�G�r���[��붸���-�ce�~�n�;����=��ѻ%�;z����V�[�_��̾��䂔16�Rك��K�l����UG.��B�m�~[i����wr�����O{�)_lU���~��ǻ��)���6�Ϋ!��m��lD�p��Xՙu-��H.��0˾�C&�������ٰc)D�����Stϗ�{+8�>�<�My��r-�Y��&*�S�>���c=>cr����$4��4�Պ~A����KI�Ξ����P8C�^9͐!����R&%�E*}�r>������֝:�i�d��3��y�Q��ɽf#Q�l��PBX��8������y�s���P�)uk�֦^�B�����X�)���g�z�Հ���`��\DW�N��=E@��o��ړQ3�4�5+��k��'���^v�h �9o���y}{J'D��ݎh��py��ȹ� /���eк]�C<[��.��ڱ]�1LԓӉrU�	"��v�@�R-k��o�.��mz�T�$�A��� g�]m �\h**/9�|h�~�ɵ�U���ȵBi�^�kr�fe0��U�pV��߶'V�C�Κ�� �SO���ͭ)�-l՜Gq}�J3N��D� g�fǫ��ɹ|єL):.-QEQW�	��Bř�}(X��~2?����,�$�����=[}��]`�!�Q�^;W��p���.��n&6}�L�\���Q�w�{y������V��d���#=�w��^F�̟*��C+��ȅ�����JT.b����u�X�Hǵf�6������j1B�L�јE��,Xk�LŬ��|Q4�kG�m���w�Ͻfo�m��%��pM����XZ�6�'��
=�ߌła������#���o0$�W:�d5$�F��ːjA��٧�O�Tx��vA��C�$2�=E�E��]�)�H(q�F��l�������1�E�b9P���vY��S$��g�Vj��|N��ӽ���Q���3C%�,�ݜD�ޮbncq����ף�z\i u���d�?d���jdS:tw�ߕ���J}Jw��n��>Z9g��?6��UBϗ�Vʹ�AU��^��N�S0q�o���\�zW+��M�#�v_�/��E��Þ>�>�X��@�j8��~S�N�8� �$�)Y�F�r\��"��ςf^J���~��o���u���sr�s�����v<Dݷ0�W�����Ҿ7]s����a9#av[�i�Q�	w��:��*ͤ����2
朠��7��r�z�Y��پ�d/0�B�����/���T���Q�Ι$Ҹ$=܇�fe��\�"�RLJ�Aym�Ӟ#�@�I(�?���JM\������J�����k�Sy��/ן�v�O�5���2��*��t�.����٤�A�o������h[����Ӭ���a�D��$��_��i#�:���K��ͥΒ�G���!n�<�D`�R�]i�C2�JK~�j��.��Ct��*��_�o'��`~Q�)��m���A�!����
��z�^���d�Uy�P���e�)����c�9VaՒ'W�uV�5S�$Y4e��.��F�a��+ҟ���P'1��#]0c��F�Nin�AQ����@}y��Į�T`!tz b�xhޤp�L�g�";��"�ipA  Za����4�V�(��@D��p����Z�r>�ʈ��U�8��K��6m6�'M6��%���G����*�z��S�koki
o[H���H��	��U�����B�u�E�&F����ޔ,Gr)q[�Q~�w��$��S��4(I�'>�l������v�Wd"+�U�����S4�f��K���F,���f�輴wN���`�fٍߞQ�	4�_r��91���*��4��D짖&������9|�'�I0�م��dc�����-�����ztx!ay;><�_~̶h��Z��w�s2�̙���-�����/U8�����H���۔����k�sj��Y�?d����~�:y�]���_�EN͈$r�L.3�k�1/�E2[�OO&%xH�"o����S�Q�����8��=��E1�Y4�Z�� G���p����I5���p�޽� R%�"���z�]�̑���[Y#�'q��jC.�&΄�P��B/=^�~�6�ǹΐ�t�]��
�Z	'�J؝��6�t�V���˚w �tQ���5��E1��eH����cu�j�IE�A�b���N5���+���D\8)(g��Q��b��o5yĪs�.h�ְ&ec{�������%M�G��
$���_�}�J֕�K���%�3�J̈ج�Cm����sU������gR��A�X�f�(��N/?4�|w��"�B��5Ձu��q��q�=؃���XT>�r"`���$�13�l�}f2�gu �r����V�1�N'޺�M����e2�Ǥ
��\b$��z�9��$ ��ۏ戈��k�uw�	X̦z �����"~jz]¹��
D��+{��ɉ=U��WL�(����c�;,��!��-��aw|&��$�u�����?d��;֍Vá����weB�����h��X~Q=?{��k	^���߽��q���1iC+ڑs���:��,�@C��/\�t�O�I�І����uh����DW�s`�^F~�L�k$+	+Пh*�of�J(_��J�8�xn�ʠU==�x1�|:���aZ�f��fb%W�9�:Z�»à��	ԑ~
i���LrwO�x��F���{<ck# ×�a����M�9�#��[��΂M��,)������=���`{ևVCL�O&�s���D�����(Ƈ��M{�m**^C=Ϧ<����׆��.PT �іN�+��q��@����c޻
=�G��=�7a s��"����4���%*^>�R��I�Yn�xk+����R����!B[��,����0�[��9,�^�>�*�a��^-�z�WPG�=�D�:�܊�S<�F����65���*eS��<�n�b[{/������p��&�
�x��J�!f�Q��Ml�(��?������W�'�P@�=���V�u��x�C
fL� p^m����F˝u��Zs6���aD뾬S X���.#&�o*�#�wP�&�.$�A���J!�]"m�f���,����枇_�;����d���0h�:����\29I-�/&-tK�<���dԌ�����P�Y�p�o��G��x����7�#�gwh��`��l���u�^T�0���(��$R�}��~���Jv�A����64�e�u����L��uC�&	�r���<�ٺU�mKu��φ\��+�d6�N;J���<���b�ñ#�� ���&������͖]@ LR��������r������ �"2��ĂV���Y�X:�RPc�ƺ4�����+�{���x��vqqI"�G��.��=�1̶��z�Y�:�� SUkv���z�U,M�L�%dj߀g3��M�h�m�y�B��v���=c��**���I�k@?:����PФM�p��R��3q��s�a$� !�a��C0� �7��V�0HW�x^}VH�����v�T�tkn��習��1���r�$���C���J��2cu:���|��
C�c���ZV��f�
ʸ~vSDc[��[םg�h���hf_���A�4`n�����k�!b95�	��`��t�N���i�l��.�J�lj�?|��м�T��E��{�-|�ӺA�,	֑���)�wI ��lE�%������һNx\�Vh��/���-��z/��RwG���[T�PR)x�5Js�e� �g]2�O�l�~lq�n�aNh�3Ot��3�g$������Z;�'A�����-[���GCN���:�����P�&��R�d�u{8�訽��~52��^gY����P�U*���)�9�H_�]�(����ɜ���R�]p��J��\�ʍ͸",k�B٪���b5(&V�� B	�Q��~�$=W5�.5��'��W���
�9���g��@��,�"$f�2'rEQ|(����R'�}��$����|9���^����%���3�5�zx���ٳ��4aL�{`(֮��-bB���U����� �bwb�����ȹ�]�TZ�z���m�-�"�#�/��ߤ�|)�9^!�i�\a
n�<}��R�F��X�����eC��Z�nM�����,���YB�fP��˛�3�h�tz`wp�V���v��AX�ErC	��A��6֮!���&B�K�=y�4 C;Q�AP�T�4����+墘F	$qq��R�"�����}���g��qn�%���n�`V'�AU���N^�"W�M���-�ŵ�+ˮ(�Cm����]�C�:Z�F��Ɠ��)3���o�BQH��3�g7��<3捼��
f�l&aA_�-�y�hda�}�WWx'@V״�h�X�,'�p>c������Fov^PY��lx�y�~_��J���I'�S���1y1X����^I�W���X{q���Wr^����7M��(\|Ԭ~!I$lԜ�L4=��u�/U��t�oi��&C���3с�Nc)�B1^�6�b1���9jV,g�҃��A�����0>4��ɣ֊��y���Aɴ�Ǣ��n�~E'(�eC)��°b��	Z��ɫ�=[{>H7�h��_b��g��{<u�S��<g�{E��|b�W�܂y��AZ^��)M��L�O�N@?�1�#�CD����������i^Z ���u�x:�>֩(�L	4���V}���S�g�W�y}��1H�
����U<ؕ��a��Zc����4��^'���lTM�ڥ��G\��q���-������ˎ��T +�'$7��:E�b�!s�7�T�A:��沾�S�|{�R�6�QJ����y�>���c�A{��f��cmu��+:m�ప�^��3�������������� ���D��g[�vy�ߎK�ע�($/�T�H,K�A���+{�/>��[���,<S4�]$>���z~�oE�͏��;q�:�"��2t��az	=����D��mC H���A#�;��rM�*�%�ǃri�F��^.��O�}*,;��-!��-k�$=z4�k(�O��ϔz�MT���^�n���nS���=���
2��'}b_ٕfs�)��CG�Md<�h�r�������-��L+mV�PY��o�#�3��~'!A����d���?�������Ѷ)��"����w)���4���F�XN�!.�} �_�1N��W��2_	��w�v�N�t�;��ՏRG�}w���!o���8A�������8��2��sr; ��[39C���Wcdi�.t~���]bm���U�7*��Z)-���dT�U�TCi��ӱ.�K���<�lv �t<��+Fl�˲�e5�Rlro�l���,˒9�����T0>_!�>Gejx`l�1��=��~u���TU栗���e�Q�_�vj_-�[���K��G��#!/�C�c�3�1jJEf�N%^$^�i�o	d�� ����Q4����$�L�Z�/]lK9mM��.�^>"%������	wfX�> ���l9�/�,@z;�4�p�{�;��c�Gʷ$Wk@6�b_a�ߝh�,Z�xu�8C��Z�t����4='��ɦ���P�r.!Z���D��מ��ֺ�'.CU�P�:���|k�4Xg��6c!��<��[O��P8���}�����3^��@���0s����*��l��NX!�*�c�y\��kT�`1��&�ۄ�N ���ǅ���R�: ��jih,�$vn���l�f�8�L<u��WJ�E�LgB�	�2��-?��f�Nx���8�M�:���d���%����ԈU	z7v�3�1�$�E�RHN�3�%9_��f��@�%%��c�[�U�2����qv�0譖4�;Y�<�|�	�J�5;��J��4��&�uz����3����*f�e ��o}�2!<�MB��%[�кX�� ��=���א��ۚ�x���'�m(�����-8������'2���J�]AK5�����"�wI�\��5yg���33��`�kA�!�3� �A��W�n���D*�����������Eݸ]���7�m�k�w��{нTh�X�
OZ7;�DQ߱.�M%C�ڌ�B��W�-����=�=�`���n*��I��V+7xE/��b"�����~@B0���4I�Ѿvy����J	bJ(�`G������6x+ߐ�'ZY��t5O��KIM.CO�0~xT��6`�G�� ���(���r0�j�γ��hXM�챙,�������l��Ыr���?�[ȥ���$*�5<� &e�d��N�;|Zm`�^e�.sY���u�<�\�oq>����ֶ/w��_k#뱩F�C��J~�
ϟ�;�T����P��=#��,txsVw�/�Z�I 	FӬ�^x������=;>���_�qsNPypV{���F��8�Z��%*�����V��MR��&:�.���u�`��0]8F�8�f�K���ɤ]������Vz	��C��计�O)j@#)L�rl��)-���H
�����c��S4�#!��E�9�&�"_Q��©��>�1Qˎ�eI ����W�p+Q�GH�CB�3N2(~�%��|]Ū��>��=�i�����I\�0H��3;M�0��X�(��m��R��J�I��4�r�� �ӊ;����L7�	���!��awpK?�X@"IR�9��"�p��+�i� �2����8 ��j�҉��yWC�MA�K^|r�|�LIh������Ln�^/�?(Q��e��T�!��%�ۄ����� �D�����{�a��k/��H�h�Xp
�sH��5(������ɇkW�G���~�2�w<R��y2}i�w��Ϩ.���R��L�$*j���P��N�m�N�F*����w"$�߯��D� �I��6��~�4�D,��6�̱��91#{y��H��O*c��Vx�71��N�*@�:̏��$��P����l�l�
^�� x.E�7ڛdsr�\跱?�煱�����PB�2,�N���aE���NKӫyj0T7m�W�!S��<r�'���S�ۄ8U7
+�Qϰ��Q��/|`I�&���_X�34�p��`d0�*+�A�y@��@��eX��#��r�[��Ac��+{� �[b?\��v/�ʌ�#�\�Yh����V�s���ܑBYV-�]Q6�6��u��Y[W�<�k��zM5h��݀�$���\���R���`�߸E	�.������	8�5�02)�;��!b�4�c#�'Q��?����d���a�m�omS����-Ͼ44=�*>���tHyM�=x�L��_�y�2ߙ�%"�c�{���K[��2����C�tv�C��:��٨���@u�Q�ARH�*Fy��j�>�B]p:%c����	igr�����Uf�^	����v�2�97�ɓ�7�Fe5�Xu�;��	J�u��1�^���d�xR�)�p#�گ��	wEpl<H��?�� ���,Bm�\�̟9�?eŗ@���c�<'ٱ:)�F�-X6ǀk{��kxӰP��j�p7�j�V�vL}n���.3�\��}U��*����h*�xa�8��Y����Ke�/�`L����U�;�����T�;���U�<��,sؙV%�oϠ�U���7�7�FR�i;~ތ*��W�-=���Q`@�,��̔�����y�w�(����b�JÍ�>�N�\��s?fc�ld�.)
��E�<'�C�����*��fɹ�����a�`GGW���uчC�vڻGp�/E��^�iA�5}�l�'�k�prpa��ދ6W�!��mv���gpp'E�Q()��?7j�X�_�s���N#d�m[���bhٺ�Φ;�J{ȍom鏑c���܀.K�{��&�� ���;yI�F���cV5O3��������k��Ra&�q�(����S�zx��45��bM��6��vI����/����bq� .M�am�<kk4/F@^�Gߣ�u�7��6t�b����[� *�>�h@7���}�ͭ9��Iʛ�6M/Y�k3���'SG�S����p�~ۓ"�5�5�b�Uj���3
Q�*��~g?R��6�D3H��Uv� �JIh��y7@o"Y�G@utg^�K�\'Y�ü����i,�BG�W1[���Q"57�$P�^�OC��=�p�<�5��`iz�a:�U�8����v�H�*YҪ��b
�L�[Ǜ�?@AP#�x�㮐���O�Ia�V`����C�MY����U�7��ߔ]�LH�k�͖�H��3���ԉ"��H'�N+�P����"�}3xLjJ��:����b̹��sdn<�}��։4���dp;�l��֨ߢ�����G��,:	�d�4��΅��OUt�J�y�~��X����e��M�X�a4�,�KK)�M���;h>6,�O�p�j���I�8.� �\��ųT5�0|S7�mگJ��S�<y�OB ��Ӟ/�U�w�"G_�zg�v��B��Ts���x�)�#�t��TZ��#���������|qs`�9�.�W�0b�x��f4&��̨�Ąt��, �p��2e�����:��i5.�񭿰0U�MFԥ����E���C�hVL���<-����K�~P���p=���:tb�p�2^��N�ݲ�����M�� ���\c��<b�B�+��o�(�����v�lb6��
4H5�1]�$4�a��~�<F�=$Lfup�W��,���+wA�3�c��No`~���(�EX/�.؆��H���1���)�ŹU��O�]4@Z�>a����VomJ�=xҔ��w�`�LMM�t�G����i���kfiS�F�)�NC��c��j8�7��SF�ŉ�_��9fD���Wy� T�4���M�+]Q:�(�9HR���溉�M�|4+���B�pL4������Λ��u
��#�q�3OD7{@4����� ˤy�bЋ���N5�!)�?}
��f��ؑ�Q^>xԇ�6Ds���Ө�;���y�����W7�ƚ#��Ț9�f\Z�E=!��1����;S�O��u�58Z�׺�jvxڃ=�ah�e�|K@{��4��9O�S�ҁ���l�y���^*+}HD��BVˮ�/vUg��{�^���Zp*������}X��êŜ�A�\�Ձ�g�Ҝ�M4�%�̴�f�5=�vҭ�l�����L�RSt��r���#��;�a�8FM���;1�� x��d}˓�����m[=��Y�n����BcL��������?�~�N$E�Jp���8�Ӷkz:'j�i�d	B�;8�2�T�%{��������z?	���ңWP��ե��z_��1֢���4~��!O�*k�>&�]�
��S�W�߇.���&T�O��V���*��ie`��v�����`��f�H��<C!N�_i�������/4aY~�k"�IT*>�Â��4����S�U*݆�o� ���B��"��Y��=}�Odîn�߯���we?Wy�c��Q��ٔj����[��ݣ.X5G�<��r"�PlwJhym�e��&g�Z��๓��'�I�������|�4쒳�ݞ�d��P���u�3�Q|h�5����}��x�e���.g8��;���)E����@9�W�}"�X4A�c]���d���������^x&��1Єe(|P���� S�R������C�o�îpm�Z�fY�>y�P����gkYߏ=s:I�bD����U���\�.�����n*=UW]iE��䖩6~̆w->UV�A�I�����;d���C���'��3&�n,��/��p* '^��P�g4�2��˫����i�JS8OE���ذ&���tr��Ӹ�$����� 1���l5��d�LWI�+�Kv����	O	�x�qw.U;A4�$)��]�H� I3\_߯K��b_�I>�gfV���W�M�ݧ4�Te^�E��r�%�\XW�y�l��9���rwy%&�w%���IH9ԛD�o�5�b�E������4�0R��k��@2�D�i�e�QW�@b�{���PopxyP�O�^N..R'1�A�0��ߤ�-Ip�ؐ6�K�\2W�L�<���[e��$0|Ȉ�e_Y��hб�B%s��^�~>Pc�3�9�ڈj!z	ȃ2R��;,�nsd�u���*H��%�닒j��0S���/��"����z :�)�j���^�a'|X��.?�Aǫb��o���n��Dp�X����f�|��e��d�Z�t8�˷�<�"�$3=(�|՗|�[b7�j�:�	��ՓѤ�F�n�P�+9��Z}��Q��� ����t6)C6�^�����+�(1�I��+Z[�(�T�DD8�J�1"�t�}h#~y�M{���=��A����SbW���t�/��G�cc�Ƀ��=Iӷ��+�|Iu�1��v>���x����|>�J��o�t�1�ϩ,�c�3�>TԻ!<�A�YL��Ѵ�+Lț��K�@L�#
 ����2vZ`m�.�O�����.!=�wJ��k��BƜx�J�k#�z�U��m���mۺ.( ����,`n�Pa9w���pa��l�j�RU(�5�>m/WOZtmz�����,	�+a�C|Ҽ#��\�!��q#��-Ź]>8U�Z�b�����6���t�	�%�������3��R{O��q�hB@�6l���t��Kգ��t���AZַM�pu�n��K���M�;�\�,e��'��	2���J�M��Z��1+�ȵ=�p�º��r1�;��bX����%U��uv�Ῥ�"���us5%�B�%�|JZ� ��:N�I���T�+"<n[X������_�ケ�Z��Uy�5��FB]n�I��V���1	o�����@E�<���S�䇙�Z��ҞA�M��1C�+D޺��z �뻉Kn���@m�)��K(+��2��1��ň��2d��t���"��[C9Y��h�R݀�pɤ>p.����#S�y@�$�/�������A4�g�}9�|��#>��1zSY��<J��,�6X�j��`Rã�֬�}�;Gf%�[�
��Ờ��8�,<�� ���7:�[L�����sAn1ӷ
�@V5	�GŔ�!_D&�N�6d	�H�P�}���iwͱO`V��c����ói̗�6�(0f���������5�`���u&^3 ���IPàh����x�*��&+� ��z�e����D�tKE�ɢ���S/VWLk��}�}l^U�c��:_�ݰ�櫆N�Kb���iVYi��\�羿X��j�\�hhu���-�M���=�!Z:&=�Ёh"�7�0��ð�2jT�#�p_MU?��D�m+w3~vNn0��p�xU� cܽX�VY�Θ+y�Z�C�|�~� !��a��&>Tc}�iY���YPե�d�-ճ�I}��rf��"����电V1�� @J^�!�B�}B����36�2���� .��:�jR��r�a������BߦR���%���q�s����Ↄ65��TF��Gs�u��!Ɗ,g��Ψo{�B"]�,	�X�#���g-��l��!�cOQ�H������Z3u$O�ڗe��#�����w2�R��f>`T���m��v�TT�ƈ9�kW�*ay�m��*��Lb�RFUj����S$��4M��j������^�2�����3�bz�4n��S�J=.0Z���C��_e�P�H� ��<Y������:e�m��.������p2��z�3��I��^�I��z��ʦx�7I�E���N�r:�|�㦒�ƏȽ ]�6����+�ۇT*���WA��	�TnVpL�@6\�s5�O��N(��O� �09v���_-�	11�.B"�X��Ĕ@O��f�-)0e�ch�}��O�s�#	>���M�9SΧ�b�ߒ_�chЙ�7�f��;q"�z�Tk�4]��k4z��}��2�iҤ����Tg	�en'j\�)��`�s�|@lZ}G�Y
����w	d|=vD���;���%9�ff9�a6Y rC̬����$�/���X�"�Q�x�%5|���F����1]-�,��G릑C=��-���FK8D�' T�1h���1�g���ey����ih���և�>�C�a��G��\�+��<@"i`���%w3���C�S ����41�������m�����Z^61�j[� �ʸz��(J���¿U6U�塘�d��l�"qr�S����\rH��a���	?���R�
A���V7�s^�����v'Ġ��-Z,�y�y��mxu�0fޥvN>��7<���������G-�w���Ӝf`��nל~�o�e [�_��eO��8�z���q��c�?���i��@��ʇ��Ps��tN������e��H�3�F_����t�#u<�Xfʸ�b,J�'�/��;�����GxRޅj��B�����*�@���g��?�A�>����e�� �F[́ٱ�q�埭�`Lb02�V�����k~�)�=���}Q�ds��J�x���Q��*O�0�}�؇4�?p>�A;dr9s�:8�~�r�b�vF��B<Ѻ����	���-��'�^ r��5�)��M�M�T����C��������Qu ��X���T�Q�a��I���lŇ�I�0��qY-��v�ߤh��
ۣ#]P�8�"�IQ'^�Y&��P�,��w�)$am�x���u�"�!\Զ��o������(Q^�]o���hY���� �̗nL��QO���vj�y���$�6D�Q �I����P�Ę�%Z:K��U4)���7��5y3�ʸ{��q����������RXJ�[�NM�wRݶ� c�e�&=]�+�^,ιL�4�� �>8����J�vb�M kE l'T`��� ��$"Gΰ�QWo�(�H4c�3��<�B��ЯvLk\�/��z��h<<�_��(���ZhX�3(�����$�l�7�W9kd���0{�Ƨi����Bz�hvT��|�-�����B�P
���e�P�j������z��?YT��_gXz7���u���_�tK{u�ؙl�LU�vAc��U�+��1�_4z��_{���������׹��.�۾YnX?���;�_9t����Pբ2��FS,.���U�/��Djw��b�I����3����s���d�-�u��6n/YϽ���6�r�5����%]�i��GyfE�9��2�*�0�O��[��a�;��|����L+-*��)��Ws�3�h]��/2�5ߝ������e���r"Ls�������)�/N��� G��4�N�ȴ�f�����������27u��Q=|o˚���wۨu��Q�@�x�޸�W �I�cbL)|�T]�fD��a���-�+4��S��ꚤ���C)����Ue���hJea��Nd���;A�q��z�V��ˈ�$�eװ���D,��D@�L�9"X�HpY�XC��/06r�2)�7yIÑ��F�a2�G��cW
����|��gy�����iؿYa���wh����@ޢ�x�R�~ǒC�n��TDSEQ�������);�:�-�"w���(V�V��$N��ΚHYk�^}�����M�k��#j3;(Ѝ���������Fc��W����d�"����n��y�]7�?@��CN��mI��f����X����d��[�����	fZf�-�h���iW��H�h����Aи�t�۝����n���1�t����I�P܋k���W;H�A�Ι�P�2�wR�L�V~�Xw3�٘��?@�9�ߛ�$(���j ��YjIZX����#���̝����x�Ȕ������J��bEs*����-j݀��%;���� sD�1 D��t�E�y.AwB���1ۉ�A�wU��! ?�н�)�A��#4@�*�cg�V��X�C�׷I� H�hJ���G%�v���wB�
9[�|kl��ſ8i�)�@%�X���}���ejVl=��)���7V��9�A�A�I[���YS��#��{#����/�o.�6��Q���b��7<q�H�1g��BO���2+9�V8����t�F��2���};���3۶��H��؈2�����S��,�n\4+�)*����{��C�]w;�4�l��X�Lf��yg%���祡e7ѿf�tp�k�M�1;u��mK��Y��Z3����j�l�ׁ%�]�.< ��C��wQ