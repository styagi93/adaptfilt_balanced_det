// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Xp8tu3Dn+V4LiezpF2pMPVFahtID5B2QmXZQdj5fFk2WEemsM8e++ZSi9t7NSIhs
3azElJqTyUO6tyt2LCdR9OI1pCb34K9qOw/Oq9bGJY4hl21GB3t71ocm1g2Im/M8
FVSuLKDURqHi0M/KLtHjkW+nk1AGE8gDC4XdAzWyZYM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22928)
bpor9Vj99/oX5MEGQpzw+Uiw1D4oX8v9ceQUa2mvY5+JZIaOj+LO9pJILBZc3hE8
Ca1XMuV/p6+VkeHohf3efCbtCsz0QNlWmi9/H2dSMZ/ImNrH7sEgpteH7T0PzmAE
fyxgZ/Gsw83bLJOfxr8ZrUMHToCnZEj6d0cbRz/9NzLnWKmu4jzUHHDEoJHEznOf
ASfczfj3L2/udarYmuXqP4rqvhcyb7qfpw83Xbp6BQTJ1AlkDlM1+hmADjLxxXOU
ydC0cgbEqrnNYF8nMo0OBDtRV9mE026l27V10OFw7gB4Bk7voW3a+jZ9Uvn2XAvW
RhFDKeCI36S134Q3dPIjG8yxCmu+Xd2cM9dUTMBMYxCha1zW5gweCr/fGRiS2i1t
V9cxEEh4vEBt4PFODVRwDbdVLhKdSOvnbTxqcDYugwI5ePnM/PK1yMYq4rL86ghY
JDOMF6EZoCQYR0ohX5wOipMNY4jGaEyxKO0L22SDomK/gBXdU4N7FCTaB8QTrVEm
wszHUSEBu+khMRk7O3cvZGjLPuwHYpvs7NR06unylpVdHuyYpIMc21zj8KJM6evx
dKZo8HX7aol/wLbBGB5/iRWPeM/2LH/jII/b7V9yNy9f3XjqqOZ/VEH2yzE9Jjkg
7zVukW1AOXU7GoqaGmAUCVByqjNRfUDmHA+G/8er73oebmveIrw0Gevvbxj48C0K
NL+P5EIP3jQub9Eb+vn4YwKR/8M7oP1OFKIZKrmJt6GAiVp5Wtu6pEv9M3tODpKO
V3mcRMfT75yX6DKBhtU60Tm97GnlzZVJxGWobnelTUOlP+3LP3hYm4JrytYDiIOf
fLyyQzMqC6waGjJfHDFWh/5rdmKy3p3Tco+K/WU6e4RLUKzvlnluLTnwZSPhqIN7
B4QLbroDs1LQ9IjOmMhXpd+Wg8/6sYZRX5pkUDxhxa6eO9woIbwpIqGHd5OwF1jw
+E8aa/SWiHw4uLH42ZekY/HjCARubSQ5kjN/v+tNqPyqs1nGTfFrTnccTsZGk4vq
y/7mM6/81ec+NWEZ/SZLq7pHT08UlJX9Y3VYsBjjfC2RjSSYFl4rMRqy5OMK1a0O
hgLaFV8lGx/Dnm22smWe20W413q5GFAjuKfwTRw38gPIMydiJxu8X48xzYMcH1EF
MhfV1w2xLcGMtwmExP5gExTSP4hZ5BW6OKeJjifawJMCz54lNqRj3Y9R88r2eEkg
vBenMiLl2XwhE1BR5B0vyT95Ui/N1nAbL6TCd+sZ5GctgRwBd40er+gW0c3nNzt5
V9iICpjmmsmzS86+PjqoGU/WfWocXuki4s7kvwGjUFvjfK5jM47AkbFm8etsE3f5
XlcAR20CA1W0BOcBl/CfrziDveq4vUsRXaMABJfXhHAJ7ewuKrH/+Q2JYI4tIYAF
U1/3ZN3NWpj2aj0TKnSUkvw9gkWoNTMEi9kFmgXmElqR14pf/1bxiChR2OsfiHCa
SU7LVeGD5UPHHDpL7QYczs6K+2vhrDNGSsnNM0k51584fj5TWDN2gLr3/FpPjZ8q
9XfodcTomC0bvbUrzFL7PSRH+PmRVivtdkw+74H+rbL0IVxL2XF5/qXkjTCpKXFo
VcAbsMJc7VStx0ALtbeypHZ1yOKL1VX13eqgtD6RJ8H501g1ist7gY4tzjbt/Xmg
l/c13n06q2zgw2vL/8GVd6oiOviJiEKLHW2IVxsDZRJJpdXRMBIZfv2ood5EC2Iu
bBmtls80rJ2d36+iVSlpkZj9d0G3yh5qS4RsPPG8BCQ8zhACFOlJLvddm+wfQQFT
c79H50kthBvBtFpCbNUF3neMXsaiJI9BXDM/JR6igSDGqwx3QQYexpxLqabUXMvo
9PXj72E8wIhI8sh0NeXmx0f6Mq8uaqiwBBEdtUsJpEUgka/7dGWtWf5QeHlwPB64
2VE6A4jOmIYPEgScLoq9CxiS8rbFmjvweuerpZSc61v8smjqgjcnhU/qSt9q1kH0
pZTxNbTy/vzj+d0Z66EZai1vDVE44yXeBxM9hZSci5vDoF4ueUVcmsc5GPl1odBP
QOHb2M+Y0g9iFyNpBeOWw4cFapTyYj5v2x208QC5l8yy063ujbw6BwAHrvBbgyTL
QJCpwJEQfQQVUjzvKJXQtgWj99z3U/DwpYjxEBpFwD1Wjs9MQ5Cidm8rysycN46H
NHIBgfUciRu+vWpQ+oGF43ZjLjkV85eeMagsLwuqmIfk0CC+AfwAXKVm+K+Wsc5K
K8a1RUsrW92ebHLdJ/CwGFjH3GNOZ8+g4/z8FHHh/Fa8LpDiJXPQ2hBBbNPlkIcN
RCY6WsJHQjRqyf6iIHKyAAGieRdMh1sGxq9zq+XT92nL0KHLYp6/czH7xHjuoBlH
sIfGW8U924+5pqt6lCY2IkOm4LsATXeZmeM8+Xiitm6vZMBPDOEO2BRiqtMgfjtD
liU7NfBNGWwCc7AbjshkASBgxLZnbH62ab2hgUW9hwfkkqZ7qpMK3fND27CYOHt/
eemqjZeSURGVfLIlb65T6iG7TvA4fGrPhsksUzI9RBqMISXwytuT7NSy67GNgIyb
Ejcw0qCge1QhE0YvBLuTSt1aD7qoOcgal8NPM10hiX9dLgysYAb8k967r+8QuKjc
9/sJR4D1Wrdd+ebojoLFR9YV8ixJ6QvP0RoNp5ndK5nEuTIbSYsI6DLwBVtApoEQ
FfnyHdQYLFIyGL6wKfjdPv9vMkpp2yc086N1iLHZlCl5crfP3cvaLBQ4BMZOTIrO
dU9t7jf1S/S2You5IuoR1XOXZej9lXPdTMyiJR5pop6i2192JUalRQnS02zgtMEj
8d9HpgxDEhq498Clpj4kh+SRLoud9JmtQn6hjNiruefg/yY43i2flrnd4WN2cAOx
M4oBNEjZ1Xh6gcHrG7kSjqqAIeEdNMdfW3iL7MdFL9o1uDjaZNLFkSC+XLAaYgh6
iWKHCV3wbrF+wecaPVHEuvh2KaIzqOvfEHEGxtbdY8SAGxetcrdzTl98A0gj8IK3
3d1JMgcaSxhByuCjbKb7v+NWMAfI06GcbOPnVQiTHAhgXv4tFfiKc1WaULMPR5C7
LdwbhlsxnPb/DauUvEc6Wj+rBpIsvgmO3N/pgPMi1Po82wYeyY/k791gBhpc0+ie
pgM8ExA4tPS7GrPadk4c+oUFphDlgBUl9xcgqHEae/3juRhT5rvAA0/wAE+ie9aA
/KBHlUtBOm4MiSs8vDIlJ47SAPj3BFi5EdNo00LZSWsUrGMHyFbhqVFcxt50pZz8
wKmTgeeESZ0RlaJscawOHzMgUtkFvw3S24huUSgMmacqqBoRo0oTKR7VztVcp9+d
d89yf/IIz28c/F5X8frL3isSKsHfN1x82OtactPQWFkf4yAgd3gRJ/Wj8wYTXPnb
dLKbwMGhlbDRyq/226BoPWYOe28AyAF/hoyF4uJ6gihsHhfH5IwURv+9ldTb5UP6
R1/WtKkr9bYiLl7xAOXBiR8y4O333U0jkCxQCzJeL1i53GXradsGc2ExKWVETlP7
LjyeRL4BROcbosnC+TsH/ORZpKb9lis/RAytzyXOXfKGNZTEFxh+SE6h760zxqv1
pWJesCp7idbnJ9kH4MTSXup8e00pnq/dKsoqkqqmSyZaY/FLW8CqGN6vN5rYewZQ
eM4rvuLdygYnArWdVVuELiFwGTlf6tnGs+u+AxqNDD1xbmgHigyJYgvH72MnkbE1
rjxIIoNBRSTlJjBuikk6xwQiPr6PPNl07K1DlDhhsL9RvmOjXDaJROuBtqGIzciB
9RS9SAEkOvkM23RPR7tigrwaxGBOzOi5g4zbwgEvYt7XAMR5BwNgap2oALHd2nBS
ThK4jdfbDYqbX/X/AVbUd4AerfcYGjaRBLqQXynA0cLzwLarK0KDX95ov1N8sTES
0P/0NvfUsS2MmyMgnOEGZ4KBR9fy2TpHC/UyStvwrrD99P++aPfS/Jb7y5F3I0XI
J9SZGJe3E4a/O4yrGXfKr0m+r2Nsidm3AxfjUiopI/KOPd0wvtr1JFvH9AUY414q
hPp4rJI5cJkATiz2CNhoKWYiAPkXnNma+AlyQnfzS9ASFxkL5dzaDYD4UWgIwty5
/cUkLlA8Zn3F+gpN4J+ky5vdquzMxRg611VZ3bAimts6fZMKH6f521mfe32oITUm
RW/pOnff5EHk22HLfftCx9QTKi4A7Me0nvdKM5tdT/cgIBnKHMtMnnpwDX2/YK7d
A98iPuH4l6snuOy4TMdwecsLIbTc3SVUd22zBshG1+WuezLNO2d4iw/y+At5qQpz
PJ4bJEbUCzJx5DG56MO+3iQa2dVP3YEm8wg35v99kbZIvOo2M3b8ymLo5E8bvTZv
n8VTOmZJeHRwn00pEksy8QG6URk9V3aNW8Z4oTGU7U7mBftr9pUslFRnVP5F9leU
3t3IvtNCCsmOq5g2brHU1z7YQHzPO/KFOg7RztVxvAXfaGwmdStdbj1HaqVDQiQB
aCCsYpJbv9CGLtp6URU+4mWv4pD7EU5TPjxn++ApooyvziMsOl8AI32aVgMSSOAr
/77uuaWyoL+HEIqr4Zl6dGa5aRU4EVh914sZoJxGYpTK1nZqyZV3kGdBb2ipVJtX
sXzCQPU9tjDUtm4UIBZfR7eMVO+8Ha6EawcLMcCUyUbyos76/bA2S9lJMX0yWyI9
Y9rrv/POZPVC8Fh8a1YUfnB6I4enVhmz3a/1Gyskd2tqaea0yPc62qy8yeec+sMp
SXTmBE+jeSDhUMI6w74fNhlzS0br559U1MMXr/vz5D6simradRywZ1UjUYcKVvE/
fWziXBV/gpPd23Dt+mpEV5BWjphNGagK5pIXwB/7uLIsc9xu8ofVaJGdCLKYkOc6
p84nXmHHN2sDj6UmJ6FigGWNbpBiZSNDoNoaGQfBUyKSaclQx84WNmEvD51G3uEB
kNok4AnOC49zFdrxi5COlJn8SDkQH1C85RFdZhfz99kjF6fw/bQTeTtzXcEPKFrC
rS/8tzgjzNb/y5uU2AmvsyRr7XNU16hvQZ3urIlFjE5U9uQ2g2xzRAB1wh0f/4Xz
7hxbK0tT2U1kEIlFKXRnUYYVuMyQATihF0NfatLrVH74j6JuZ49GXIbRRQ9liZ/b
Bw2n4wvRq/6J6IdtLgnH116dN7+Nxw3GzVmbvmPY0fB5/C/bNGu6GExlLSiBPfee
hwfGV1Ce3W9yroiDCDQDasRXdRsH9XcOUnnjNmJRYCMJZXxbEzLGp4ve6eyo8NfY
n98iP+L5tKlU4tvqoo0dmqTFN+YX0QL753CYKcP7lhRJJzXxAeaVXfV36VnUspjY
J0pJWAZDMZRdZpJMTzwkoUIUvBSGJKNwPzO1UHgS3q6Y3r0fvStm1a69qR6U0z8Z
iyS95juNRXu2eUsqd1GbQbHg7Uoy+W0WEGp2nFeSmvzr8KNHmPUIDBVk79biohoG
9CcxpwvsC6Tj//n4NgDkBwZ6nKeKCAnLnd6kLJA/khagW7a65f4OLgwEeUoJMFAJ
RImfybES0zh7xc33TacnmDFOnZbb8BJs3SO2kShXK3E1jk2px7QsoZaS5ug8xeps
xS9AHPhG+sCVLpU35NTbxudA64QGDyr1LHuNSA060lEl635Omf98UNSKt2yfZTed
yhB2YL/IjJcF45r8vxKsQRl+XJXklDYdiTJGhE+6CEFMWGvqx44kH0RiV2JmG1kd
9UqPhAOeQHRCL9XjInD2EtYtf3kxXWnQrg45orABNcRynlpwFkymqRgj7xlNx2Qr
jwSPvWJ27na5Up772hxWArRjDodjldLZsM6MUxrrAzfU1nIFeRC6NWGzqMuoLoxl
sUQZbL83LuhLjqZeMc8HrpkUPuz64gYsGS7u5yU5G804mTfYDBnzQ53Y3dvo+f23
ZbdUpHCvuF5eZT0upuPVa1D+StZ7UDXrjZFdz1N7ObNvKV2ptLOlisGpUxTSfLU/
2UDhR3yS9t5Lpf4EO25/wNVKEC4usDqgpDPglg3IBcDIXjeXfNz3T1Gx2oDXA4EY
DoA+E928FdFAG2P6AfFTV05p+Bnjrpv8p+r5zNQEoGLLW8XhSjaYpcAHJ+n/327l
kq6iVaLkpZxIyrhG6B1UtW7Vu2hKjvilt6jKFWMwL1GnLCaq82g3McGDQ6AIByxB
tyZTLAX5fQHBGi12qygsC/G2cl0VjTW84yIKX6DwpaxSssPTxXA19ZLuk7fBdmaz
XZoKWAlom6XeVCAKH492XOpLx+RMlAPtOCLUFcVVVxZha7roXLSMIlTHA4QxSwUK
qEz/C14wqmkMzJr0IWu0OnF/+xcbvGVOnWy7JDKVMVN70z0N1+tbyp+Bx2+XcR/r
xyhQP9cK5FVc1IAqUt5zudlzUFSh7ENmtJKtJJl1pPOYwlNj2Zze7SscJy5aAZRA
qczO3VU4eD1XELrh3TNmxHyzYijpLb1RV0o7yl/QqI4Snn6e+mkJpYN4iJeKhO/4
FSXP46lt6xiAiMytONqnbT+C4v9jmoZ2Y5KSPRQPjA7BsoHiA7X4EZ+z7Gsbqydl
59rLnOjqXQTS+i0kG4w27uHhY/g27jfWyDAIi6m6C7ZxEyi9yT6W+/8yuH/0RLUU
UrScCxr2zbPSrO/yIPl93NQY8K/81MLSBtm0Nm4lh1q5BpGuaxfl1vSsHJLP79eB
6X+vYmNWgXFw4bm5e2NH1Zsgy1nOmRBQa/WvQYLBsMUWWCZiokztbeYdxwGSbANe
eOTymLXSymfk7Aeh8RjDUwkPRmgF0DgkDZ1xoYFuC5fOVfjLWN9vSvjGG1gctwLV
eH3yYCP6Q1pnQjQJjU1PhMeuwS60Sr7pohVLJAzy+L4qp0vNNYdOyse+m0/7rCDq
bC+R4osQDILQqJi4emRYYo6QUJWv+o3TlCujvJrQ+4ikm+Hig2gh/6gkCQtwD+r8
+g9DglEDCqsJRVfNYittT4z2qMAnSFY9wJiowTqDA3CtKj6v+UPA6eTgI4MhhViN
aBduRykRKCrSuTjbCikGdGqSB2DSfhcUCj/X4WfJYAnviVJlMgNkilicWDKUn6B5
5II0NT8E3BGRN1al5xv6ROdWgO2/gS8PAYWMLqFX4DeNtoXFet4qIdKrviLb7EuR
1j7m8XUoa9A2+EX4LGDzRiw7wgt6iJ7uxceAyePmkLIq6G3MYATQv9hQvDkNtgKT
Zd8kR9E2eMUQGgem+NNfvrhIuoUJH7d4deZcXfukk8yFgNAmjEVOcwC3uNyzl3sa
gFFZJW/FxO4fTa0LEgPlwicpbeJOGPq4/UJ3cQTqZ5C5Lgz+olkN+crnS79kxG5G
jLyXoqThJOFvB7mA2GX/bm9RTK7AaNlhbtgLB5VILsIaad/WBEmJ0uOwmu5bgdMS
1rP6+B5qanFf/fd8BN33/SPgvhaC8lL21OqkCZUfn5/GAVjXjsZd0Iqg8OfEkeAR
Oxcrbg8LzBFyv8yHrU9GcpFQiQyDxOnORJs6iBz1G/1jEBxJptfonIFh366FKAZH
Nqch7KQiX/gRoXzcg5jCZ7k4rS7gVJank70lHMi6kjI8kmAaz+ErNlm9s1dpd6xe
YmYPDrEbh7df36N3tciRVyecqpVo964RhdP2LmSVaxdfZIdQvWzEB647tZ5KEWPF
8/gqPtBMvmisGEbdhFUBrWpEcVPoxyQNX6K0J4PAKwTjWTUhMfVHxMVZV3Xb/0uT
NyHXWhQT4Xw7hzxto+3fTfiKzjcCLKpPf9voapAfxxfe6UC7lHAVvvUFyt4v39ag
bD/dLiJEUK4+LpmLtuipjugF6rvRybx2eSaEV8BQHwW5nwwMAONexZ44Ne+DlJcT
4AAavC3fvoPVKOEWGbmVeBB03uncQz8JKeqtdwtbDlsQL0Z9zkAiJFUAODZ4tqVr
aElFxhf+IrmSXKjGVkkxZ9eqZ8lTpt7glHcTm0RY1VOHAfIa1Iq3wqlYfXHrSa+/
R2lq6yFyNPyJ9zRUDkskS1APoHRCJtV7U9Qf1pxLxASbzW40O8Brpt0ksIAza0Jg
YgFVTEVNFQYrXMeOfB5XUYdvglK5O0W+4zzhxq6a2ikqZYQzBth7Q3tYXzT7Qenr
6IVQR6ERenpqiZqevPWNyCpkf/Nqx/vhP9RyPbsoBt4r97maBcHCGnbXXoYI46HP
09ZZTEiPMbFMFJU8AfX4GfLKkEVh+NZABJGnJyKann4x3qDSltXoZ8N8Fij5+kat
YNTe1y6wMkWdgrtCIHVtcl+rl4oimUeCWm7fHLiLofI20W3ACWqPrii5ax+ltSq0
UGHuCC0IQhCikLDS6hvnEFZzlq90/8/TYjJ+Zf42xF5a7HT9F0+oG+4mwKnyHQeB
KxLuIj55JtADQYlKBB+ZlN6ldwRJ+2w8wH+JUgZKF0+Pe6HNzOJCsfEvfK/qrr2Q
Yvm8n/fU/JK0/VenLOAJLkvJszgEgjmwek5VTr62GQBUqPInL2mJue2y2DtfRc7E
pI/anX+iCozWDLhYO2GAdF/m8JDQBiwe/YJ3ifMKCyRrvCt5QV2SLXyjOsUsfbOC
6RrXF/Toj9F9LkgCCMgwhXds0J/Kku0EAORtGBcftI4vLJ5s4Vi/oUABa4dJlFPd
srrJxkj+dULPEbdBqjl8+s7SVfX5XaSuEBUcKDEZcHNyLrG8uuG5W/kGnv2qwySj
pHSp0H6cbamv6YRDF/LS90SiiGQqU4IMvcdrOA942yvwO2kCTgqPQpSvyGsE6n5Y
fC1XnI2OUL3+AotpYsDa9huTHjYdTQhcRl4AkZLVoAoASIXaWfqDeumzKl3gT/5c
Gppyxpk51xm6CK3iDBAo9h6WN5AHo8D1ADGYZiPSYCNMEmJCPdCJUpElPjDKdaZJ
qy5Y++okZ5bLgalS4Uh9aC/cW2rrN2reXNUUHS1tGA8ca/10r0URUP/AfboNzwTx
npCEQaLYxj+njvCJMty5jVMplLfRAEq6oPUtqmf9tiS+xjJHypMvcu6Gcg2Bm871
TEtOvlEVzJT+Fj2BoQ46XiliiI2l0c0rkmm4sDy7NcCQGKAPwHDsawm9qH9oEMwP
Q53YEAcrmUQgV6mkiUyuhgTBjwcxf52/CdAD52CmYoI2jKWu+EG9hwuoZObRzJxe
EEnXNc6FXUZG0Aq41cXA8x5weIzkc+V4wepRwPDLDfJo2Bw/JQ0GkGIaD7TBWVUC
rCLHUN3njMs7vrUhKR3qvyC2YXpbUrY/uqHir36HyfdX/+S/XwuF6CGzNfXn5pkt
w4o6aSVCEHfTfgpqkk1Vsqo+1kqUcKINI3A6q03hsVxiB8waZRnvpoMo242EsFVY
g2mHelxRAltkbJPncSwDzrtfz0Afs+/1xBy5zPX7v3el//HTBbPqrzzERlqVby8d
A3Z9NIMjGvcFbgZmGw6wDu/MUu3cCqX560rjZILa/fziPwgf0+ZwaYYEK22bUUvd
pRnW3us9Nw6LF5ktZ86A7Z8MiGkW055da9orsuT9DAS+CHOBeIP6Wp2aXy5qtx6Y
rYM7al2a9GSnjJOzmxSvIWOCjvaXmqEJ2xfnlnkKQjGnJFwdZ07fsBqjxfIjOtY2
wHSWSJaRjK6t5ymi2gj8C6fJuEEgR4afIQpmRzKfZ8J/M5Xz6hh3HjTf1kNDNA0I
XKEEISAOt72FZRq4Zltn0ipr8Do9wTrnnB/uyb6ISb6HmzJJk6/nHnPVctgp6Nmw
liDU2YSoSjXfgTyQLOTySRQMa+mzGAtJRa6VmuC1DUNQsK+UasMewEoBTuo8Z7AX
tMSLZIu+QwIy6SpfxNkIRS8Cri+mX+xRsSAq0JElPq+n9n7t7qZeQ1X/hxO+Pclz
3g7ldMPpgGIohOOfvEc8FsQmi/q2vtL1+/XgXn4s+jjaTZRDWJ96Wyy02coKY2Jt
mA+1JGbtl/eKdiKWw/Ulv7vuBhr5IN3npoq8BdnXQJc67wKEvG/rQA6AEU0BJryU
It3Ux/ycrUWxznqvaD1MxxWu56ARK5TLyYVrD8ux/SMi/+NGjp/bqTQvdWk6G+NS
wjipom90Fyp71bDiNVwLQGD7/Ox1l4aENgh7wjzyR9Y1TUkyT3NqOxm0CYqVsUOz
SdBcb03wC5A1/lSzKXYHeA56hC/3O6t3FSCuY9s1z0N7wFm3mbPRR40khU/zxfhx
Y0mNPoyr25URg6PEnK+0dsjZtJQQH+YJTaa6lCcvRXDK56JdewOMpt1b89nkYaZH
TtMS8SR12RZWJW0tBR36noumSQjlPahmeBGwo8ERofhRVEr2pZ4ZKRKzk5Q8FGXO
bdgSTzyaHODrz/togzkvQDJD083PZc4e3d+yyOSKtE5THJaWVlXSMs4LzNFX2zb1
wZXM0Wgpk+/CFVpcLwsBNSJeEm39m0VqyWnSMy2wF5Vt63kleepJiTj7Mi6tZ0Mt
Z7zGdJ5hUbLaXb2KG3Vqrqs9TYlqRDx15wDCOBSmlKvGFS7WfNHS3UuNloPrNTXg
3Xx+SgnKEKLYT8Ee9JYkLrDOP3vgbPRER9gXHH8ggBPUN55PqmkZakmP+40Sak2E
p7wyJ6rRLdQ8KyvtXReNnASGrMMhD+TIibCrXnyga/Y9nWy7TN2rDURXJFiLMMsH
v3T4r9cg/tD0gyXYZ18Wlgi/bx+GHcG+U0ZrLQWjq1lsoNywO0RgBG1nM4UrdcUr
XPQdrLvn15jBPMyg1ZakkRtzobz4zHrAJsluW3Ya0t87TsCD6G3sBMLFXiQRdhKd
4PNcAy53SGo4EDD6i/OIfIZHAIpQ6fMgz3/IAmKcAVRRQu5pIZutZhgrIeJeXP/d
HfglUAlAzA5/N3GRnnAVV3X95tXjNYWrep4uREjG9o/q5qf2cAJT/FcT63eiQ3g2
gtmlONafnUp7taTgeiO/cYRyFe8px51qrrwQTggYdc/6LPI9c9uaFZ+YA4AjThKD
T0biz/aKySnpSKcgo4eUqRFfjiob0/jfGia92awtTWnEZ4N+SYadLKu6wO8+PSaa
yeQq4czIN7Bvxdq3pnY0M0W44pG+lm28fM+SqKJe7o0O9UwmTehdM0LVdue4qQ/B
O7WRp3x668PpCStAbezFKA7xocwqsnGj3AFo7w0Ls9WrbXSI/OJYWXjcIh2KlJn0
+bxVbjHCsiQs5biwuUCCglgBVy+23cc2oUU8TFmE80+uWqbNXSHVOWmE3TXcV/Ab
djeW0M/qaSj71BXE5whkyrLgjQdA796Q7GYqAEDS2DMkA+AbwEv40wi9iwQjpysj
0HMg+n4qTTCqaVW80Y+ZYYwMAfdm61X0k6OAcfS1RlFohYd6K0fuMv+FBPskrZxm
J0N/6wUwhAg+9VHrnibm7r5PASS2IbiGcUhww1M9XyR7YlEPUnjMmH4sFvXPTIyP
U1q6mwh7tp6VaVhcKHSxHYATqhv562gPJuKA2mOPkubyKocvDqWQFc/nL4wBLRpF
HlR2tLQEnoG3TAPkdicR66LburGYsLWmBFQHZrADAo9Qkh2K7WLDxHILbDJVviZT
pXEUvNbcFgFOl8czMbFBhD2h9xbntmC6h5OTNCh51eKfCb7K0UUTs1D58cT/ZH5H
J+nifmVBI7wj2fLtEk1UfnBpL4bMS4dx0FOzVrj30WAHbms4REPRxtth99mBzdDb
P5O3FXzu+YAE3D3H4qDDqjQnjFBTQzZtlhNvg/C/h5VvKowBCGuIlLmq5FtgKMmB
yNcx7WV9gHpWxqD8GM2aeg2t6URtGDH5d9xJczeVfxK2JruIB8vQsL/0Ou3QXyyE
QjF1S9VF4cfVrqGzcOoPIa9sO6deCGbBeKr1piQ0XEpxQmgQ1G2kST6AQ/IeLv3a
ffGa+N5tbzMRkJwwPlbIhU7laJimkRHU/g9km9Ekn1BESilR+USxBRmHs8/Zcx/t
5EIXO/Zr1mOXjiH82kwlvbg+tzdrAbYopAfn+vKnRtD16PDDaeBPyxjvS2bx0nNX
y+dBuFpNX2bQBGG+mk18MceUG15uva5zBK7liwuRid64NMk6/eXA+NWV6tQ3e4e7
umlNCJyvchH/XvPSt9v+ZgSmv8JzhZNE6YSqbvBVYsazv84vlC8sym6l69Q+JtMU
lMA6u/wjVG7T29XXT3TB2xKIka28Pt0jM1YT8WbMlq0RTyUqclDvXLfAoxj5oyo0
qzv248lrJZB1r18XNxdO/pEoyHYY93aeVnyCGosTIUAYFfGxwq9RGkmgx2MGBb1v
lelw87GXlvU+DCDIa7M94RfS8ACA1PR86uoiyvb202AinucOGFOux17mFFWXbjKG
pdKNt6T/l2OIdwSFvOaVRvBv+pU5LfFbITlclKTIgjYbrrhcUkdKOViTbtTlaoD6
tXYakS4slBFUdoh2Mb6CNEItd8jfCUHUgtwKo9uNNS8/P2ZS8HNE+JRKOcHSjFkC
R/gwnEq6hVt8G+Uk0q24bFYDzblfvhNq5qznVUeM7yQKoBI3hGQ8n3Hl+fhOM4v7
moftZmKEAyFYHMSvSaagy3xBPZTnjMyTC9kHPt5xvi249MA+uxDi+Yf7coOMDH2H
f4xWhV678xnHs5RKp59EwasGRhag1yh1Rlq8u5rQKQp6g780gUemsz7t1oLfuxg9
pBg5S0vJoD0ny4LWfvkUIQwGrN0NGgFUruL2mnwNQNglqfJ8Tc20JWlGsTEYufj3
k+tnEUVSZ9D+2Oa00MXD9RsbI7i4l7mF9DOfAw/qgj7gCiPDlT+HeVWhfGBbTxbJ
4lEGRRzWPqhl0oo/vDfk6VqWoA6BkzmD1H/MtotflP57fIOt4NxbRBFtvHSUB5bg
ZYV8JOlNNM4jhALXXscmbVx1lQM08ba6g4lIm9sZ9IcY9i9cr/x62B2LF1cASsl1
0pvg3t/elZKM3jOZMsntpczC3BtzJdEIzavxOwwZbJZhwA1DldbP6m2k83zb6f1B
VM5lYHHPOIQGDPdmDF5ywmTi+ZB6oYNiGoEMf0c+mIHINmGTpKERO8b+OYnQ/VF8
T01/yUi+/rthqsku+XlbfAHtQ0KC341oKJvbZ8K3RW4LQwqK7jaht75iMgVJxDrW
r31YR2X32V+wWHQzPFCUcd+9aPJWpEjsIVypn1HDEy5JKpLaEfPf+9fR6aQIqklG
cFX07br4/OI05eVRplrmrGhmbAz12YVZOeMPgjxwZH0tGferGVBJPP96WfW3exTh
XXP9e9Vz5nAi0csGLDf/YYjRTl1L3ENo1rTuZs7okFjTAMYdnViIc8aVeXT7i9tJ
aDUQEZHJXC4+IC8+5IfePsl0K2tSj3U/7bRtOJrLKNgKbpGh/u2ksrXoM7wa+Bcr
dCmkqeyHB5UPYrKlFKUBgFHvz8ngm0EStw7wYoPosGOOUBDAJITzdJNNaoBPKT3W
ioiNtFfF+xkrufe29pAHNCxP0aSUZw0I2VV0EEcQUzgfdEkWb8KmCmYcbVnEM9NA
d1DTDgZAHb8jh37E+/0XhCnP9SWevZkEgyFApaFEfpXxf+HzNMgu9SbsNT9BWfGp
PuZuBMezHqwlnKFz173uuXko4ItukH3FBEFIr1A0Dl6WmLE//A4AmFn/UHK9qgCu
9/80/VPBeaJ8NVgKmkv+Hpc+BXacKHtLfieOjLyLESfN95jXkGsmhA3aaZbH3+ab
OiEkBDftMrbP+4sNJET5tJdCeL1EEK2XuJHtFmqMfZkrtRadUcTPRdpSqoy1Obbs
Sd4yH830bWZA+XTLGgP9dMIrAFhAhDdNJov4K4lVZcEtYKcq6udra1CEuNEsN23r
AT8MP09zxtSt+Z4VStZnptoD8xJRFQB6dV1JF5Thuy7AieUHJA3w6iP9lhrUDTVp
/kkC54IMNsavdzUNgcdHJxCW68PteZE5YWaQPMQqBgKvo/U5KeHpsiWzFDulPPqV
rCAEB6N5xIm9jyqaobBrKK30TNQ4wxX6RN3xqiMCQRJnFo5FTX/iqtSmCtct7crk
UGlwyak6EMdGcN35O7miPuSgNhKokU4GbDn1tr7TtK1OIOEIFGfoJVjtj+8ggX8U
wh5h44Qu+d04sUh1qyLWTL4ujh+CVdvUP/RUCh8Uz+JWIZzpxbn+hUCkk7YN9mw3
gHyiEgWtfWJqudxsmKe654V6Cu76+LFeeknC7xZqGaRK/GRd3+6RV9iQ4u1NG6vD
Vn3GGMm5koNDsp25rLfk4xjldC0BUhYQwnGnI/VFu1WFFFunMkYCecJcHtdi8IIv
fjlyTCvAaLpc3+PI5AfJ6hb/ytT0NAukdMcaGrQoWkLDwySG3LmDk/VKG2b5EWIy
SXcx8FlaBXHhEIlHphutLs/XTd0UgP77B34CkzXYfGiVutGemDQ4xbmLlyRlGNbe
Ou9dsf+BTAHZptePZ7JRiqZP5ofdu7EGCSTcBCbA07AVO6P2ZWcOLWJYKykDmXI2
uOOXTfyRt4p7mEVgSqsEo1qVZPth36eGpfae03N7uhUEwMLNOIfQ/oZyi7YGVDk9
CXLBBmtc524XFVgczqLpIXATuphQnD1urothFXakemqwMWfYI1WjtoRO560iNCer
jJTPHzDjRSPFAgB4ftRApZsAMId7Bytpso1KQrU3p/ALBawJa0ejw8tTFlVXYNWV
rBDFDwKqtIUlx6thfiqnpUneiTymlmmYdGdwZDJ0wpVW+nf1/ajmSJTwTxIiNK3W
6lVYr6AyjsZyTr9tq5rOWVn+hjf+ddc478rrwNTR+lkAxDaQHHlXw1CcZxJQxbyD
jz1emWxbxgWwzY59zcNAu23+2YNjxbBN4bmUm+1SNH92NGoWo4ufZYtCmwN4+Z5+
Q4ZmSz/0+vttEDEHT+k4Fd3im59pC4QzlIFqslPiNnUg5oNSJ36CK10fRvKyqaXV
ZJr340MSfsmXX9yS2ANmssjnv6nUYikeIi9QSOkFatwduujN1kwCDhMAF1qTGWcL
vwRnKepuEyDTsTQrMfhPgPZvaFY5BYgEb0zWoO/kJKE8RXbw/WdZHfVwCFGLEq1C
/G4srkUPEFvk9vQ1eZeIV29aFYOPcSgKHbt7KJ7rabF6zwqGlB1x9WvHFxaLG9Ce
u2oJ1DTMrHLxiq+8s+wJP1nB6NS5wfaTz5OlLtoGnh24DKYNOqoxatluxllmJAJv
twdBZVxVcGIT66ahlHPYWpvOCoSrV0bq9392KMhMgwV67tzwOltsHNOulO5tyF2W
rMK600oLdhbNvq/CCNdupgszIWsEVlsbsSc5jeQU5fWMQDt+uSp2KiOmCmMqqWYB
GWD7xQV/UBV3a656b/vowZLmDRmSq7TgUkFax1g4mxd6wQPBUKR2cXg87RZ29xd0
nQBAYL2fHqC/7fcUeIdNONwJC71fFJvjNVuLKfQlnAuayDzVnT1WE2BBZdkdJR+d
wDoHZGOO8YewoDhPUEvtTPcw5ByuMXsQVGk9kjtAel4K8QOV9LlLcF5U9vOOssjw
LwSGiusZu7ko8diQwcjPDK+2RfhuNU3I3yaotk/9fnn6shLxpgP5Py9UV+UNh1Q4
4UoEHbajNGiXzjp0grsuUvybRSnyhZHnjPlubE/ssCqD2eNewoZQDqkt8GwRIwUp
RuFHk3iec4Jf/iESlVwswcLUXV0hYWeOoIF7eJkdacq+KVBgIoISu8fY6AaV1n86
CknCfnN7sGhkplPql9XFE/y32qw+jf3Gabi7WFhDP8uJjVwsHtuLwbqxX0uHzYDB
ZwyD8idptMA+iil0mgP4vAREXvjTNaFyvWWuMV3KBw001PLQkJWOXy/TkPhColKB
LmouLdaFftROicxBUy31pYeskIbl1dy+PqEjeNSVx0NQ+3LPHAHmf3ByTSAxjpVG
8h3jcIwka/S6whoudqYye8XflvSMfbVg5OVODoymVWBXs4PdB5y0/NiLlDxbgfbn
G0YtXMw2dCElSa2yu5Ko2Ch3KipF1rrBiwiTqSJvHBtX5C12Px//2CwEroBM2emU
A+240nla+ilptRjO5R6SvLEu58SZ8rnVFEFP88ytuHmuIysmx+854DHJHyH48nWl
ZMS143IsXGYfDff3ij5g6+bLeKlpkUNyS8zdeggIEgS59vXWDzZ3E1oPgeNZ3S2i
uV+JTkq+Pk0E6nktglsVBCfA/Jmi1u0xArWzLns/mIHpjl3K+7LZCyTGBBMShneE
iVrsGAFya2linOMsqfaIxiPaZW6FtkOwDnfzEhMypCJTdMo/eOQZmnP5TqZ47LN8
t9Ex5ME9S0KyLX+iZMwLDC97x6I5EZLaHEDAPz8j/YuYh9qI1wFMNKz67h1ULUHh
fu4rcS8oygpMCvMaxYBJSFTsS9XGKjs6edUphPXE/3EUZaL4H4szbBgydQ07/m7D
YxmGApyyXLl+zy+ojgn13kEkdR5s57u21EISIob6nNPqmak/yYuQ47dY+AsL4dbZ
oqSCOoPVGrRY2JYu/Mntk0n7ZyqbfbfC0l999UHLoDrPCN0oiKnWxap4pOvlVZ/6
KR0r3e+065IL7BkRpiWOZqAftVduYJU2RijRvYz0z3d/4Q5ti4j9Z9mBuQweKH+X
vKgriOZYJs3Piu69BJhkhtQKUKO0/VO0XGYPGuIUYgr3r3DuEX2iJLLIgwceAPUA
VX44HaXlX8FZ+ex520yb55ZuH7UQwJ0kpCjSp6BQ3Ayy2f9bXvPoMhhbbjROpfVq
TmnC3NSjZHBp+/lXYLJPRxXMQiemQwGAAd38A8BlCc855EV43d4DlIzkf+aN6T0F
xuYJP4/92qfYmj91kY36RyINVDxCkWU6aFDRPuiaOazgvs6uyKZOsTduqOMCC3Wh
QOMftzTB3KKYBCnW5DPJubbl53JiP/XEFS0GZb1GkfKXFjefN1qEKU+1iIu9iWzm
UBZ5tLEKa9gVSbXRnVl48ANQZ5duB8VF2Z3E9LY45iH0VKGawcVLh902BbNN9tnt
C0syKzeTRF9IMifglwULg+rIN6UKKo5Ie1uL+YFM1MkkK4pMupUKIWNC5Od7to3s
TfB/sXLwJuRs4nk706oTjDFD7DFbtTDr9RYG1dMrQKLcRCRuUMP8ou/aMREl6EFe
wgT7f6tdCkRRoRxHAz/9v50U+iEAe9eYsIByNFSl2/KK+dSyd1zctxu98FwlWxV/
eVInD+hkxDpeE+qXQ4XF5XdE6lh4+5DqBPLiIKbTnRM2tCU1BIgFQ7ctOcAJU1Ub
LjhSMmJV1OO/geRv+IYJ6FWn9/FI+RGzTPtdl8g+3KoFhVK0CDWCdJjf+0IchaFy
GnH+0jpF/e3X/4lOiPFicSMt1vcM1VVOlxWHFCPhLj7LgjRYtCZooRhhQ1qKpssZ
1zA0YHpexlt5xnEOs7SnRbyTittDAI7Gf3kn21mfHePQ1f0p8+dwq8LJEMgKaKZ5
27gX4l1S2qOgqiMIa2wZ6iahfecmNwZtZ9e3dfUY2nPW41XR6RsvxZqUvbhIufZV
s06xuhFuBbAxytXXEMuAXBgFcr1FVoFw+NTg9kmTOxWp++eKVWETMVkOCMT1jQ+C
COU1+UgEYU3ISislwxvoctvqt389pVrxBtHwswAoxBsDwHJtkNAz/JZczcmPGNjI
gwA/FESOJYOG6F9Fn1pjHvL9ooEb0i5N+WeWvgJb4IEZwKZFwqBYhx8vekfqDK9F
fEJDvW8pzE/1Z0efFdpknApMuJjB5yiTPkGizCSDN405xz0NyCom+3j4Xd9ijGuq
5DXlYGVEZwxqqTGpbsuH9XXFWFMEhfjv7gmtRL17R6GdvD52Y/GcnzVpHqusMVGV
o20w39rbp74zMncAryA1kLomhXHB+j/W9/kcbRoDHw0zldUIdGfRHi2nJVwaIR+Z
zXDjXDiLyr3EC2QuT7plc8OAxFjIu+r6GLozYmaxLAIaD3BLG22zDKWV2lZ156TL
bsbvYUs/aQF8kQE6R9zCZFq+CRnlKGJLWqzIc6D0ciUe1A6+b+arj5Odj6m+H4sM
9j4reEHm1l99WY9TrG3TimfjF94JiiLxaeHiC96PM51n5hZfg7dCvCkiwqg3hMkd
bLeK3c3lddoCzq+dkuK5LegRs7S9kTYG5SvRCinIdg2WhOdiDqQbnxFMz4Qsswdz
iZCFcq5EDTb7QIk+/389inQ2j3jGzPsWmnUrfi5oVpjJUJx1jCoQqP9YpyOWRYrd
XIPFVHn+T74X9jub0JcHSSmXJ5H2rdwnW6oPbsC/BjyNauiG2n74p9kx7Y+iU1zU
3Uqertu8hD6Fg4IDnBZghe4hgMKUlWVxxf6YIJYhYvX/bTX9re45BbUBsqPGWaKj
Mvr7lp91qgJg5L+mPvR8eEQwUV9KUWtRp0HWik/DWKxrdBeNWmBxddo4IKqC13Yf
q11e20ge5JGWgdgLpO/yUCc0Iw4yu6dbbtkGk7WkdSctfClbrsOo8/iddzM4t6uY
d3xs+fYq9PDiz4BoZ9nl5qgQZf9Wfi5bHXIRBtgp7jeBvP75O/WRqmZJ0MoDpOnb
8tgLHDIIHa6/J8hXzemhPPGwQqvd7YK0JsNk4e9hHOBIsh6hWcmVPAlNAJMK6LDJ
o3L0l/9gq5e3Wzcv18pqBIlbm9teGuDslvT7fqPYBd5YRoB0aqq+b8W0qJzgYVeq
3uZ94CDlJfdDBMDJb+5gsiIEfxOL2hqKbmiGumvBjpsSB9LB1K58CxWCrNT8wlO7
tWKc93i7ahJ3gP5TOHGCT3y/dbZLdHeNo/J2umnfgEN0YosJlw/VVQk8hBBpI0uA
1glcd4Sw7aWA0rk1W3YvDeX/9G/ezbSs0xJlblpInXKGKF+2JKxwqZw0072FRrry
KegPDnTCh6dUjqeMLaRKYfmWzLNXezR4vUEdRSrHcZAekBogUiibJW8uJi7lys7t
zTMI9l+n4lnA8erTE48CZdSHXPwgfvNViKMHpeYwXkX0GENmwXO6AM4ucoaitdMy
O4qMHEmqJLu0GTRLf5mC/5ypqhujzi9f6BvKsfDcKN+CDo2jtIMgWhJYURhLAcqN
ySVU+PJI9yVFfrtQKZFg4NAKAsVGAEoVUjHhOQjsemp/TXij5+1s4Un/Oa/+M90b
luZIBo8DPHWvgs7aB6vHssaPUXH8i/CSCjc+IPv3nxvL2Mr/emWstptEtLkPzRqy
Fl/zQdxRYYC5r8a2+R966IQAGLB4jGg8Q2FW0Dac0tW2KCwokRU5iL3wnUr6ADfE
Qg55AZp7VEOnqjwFPa4x9gs5YZdNZwrXUg1Il8oWTPU6B1/kwp4P1ucTZIQPZnmT
UQamgJHOZrhGckz0BkOVLImSOIzQ3lG62SRFRcPGauOr+3EZDHlB5PfSDfE3Iv1x
Se909o18VXYk/+VCFE/k1HZwbzRV7c7OTkqC2SC10xHjbsLJtzW+Fi3LydvW/rfs
FM4wzO/M1Men6Vc6KuwbU+mB3kEwqC9nfWPpBd/Ynq9SuU7gLBigZatlV56UHMa8
TybIRohkClkshxJaplzVen9Pvjtk/uvSlz1Og8LmfJ8UTh1daXq6IvcyWj5qSFku
EMtji9HZvr6bmPdJsmjaIkciWFEQuJ1QsTWG/nHTyfbIC8BUnhv1aKHyaWDDE8Rg
FrO9ue9yLRxIJ192oK56VnM20eHcN67//AP2NgyN3zFkzT8dHqQWeK+bWLTbev44
/W6OdRl0WHQidzB6UyNrbNjvY+uRxScAW8nLxitppJChQWpO2I0/Oyzoz7fC0V9Z
bU4jZPg95UcP4p9WyHlEUIGfxPLC6Glpqe5qGHVH7A1qaQm+jFl2GEjf9t06PoBM
IbOtRCb9J/u+I+d6opQs/LRGBYXMaABGBcwXM5D5uHxWb/umxLB/qqPXKtdz2wkW
wpXZwB2mxQjGqavchiFfLpfirRTn/v+OOt1e85F2w/1MfMLSf86nQNlKlO3xdaOz
AJQ4DTS9k+kiLWfHHeO7xMlZ6/bkfHZMDnE7QWrmGL93u3Xd+ZaTiWMnRQzc6LSO
CMb6bbu67PTJhFRm4pHc0LAISjQikZdo+A4OAIg2erTcWZ2HLD94kFwjcgeCmTE4
DB39CjTQYQo4zJsDeWL22pBJjNjvukZFUionPAKXowtUE1Y0PvfBlAWD1FbwRbLl
69vtbfeVTWZNdbYzP7v4ytO/++pNaSsZYgyY1piWOlugsxi9eCqasdrLdXHhlhaW
26GVF5IRpuW75+YoZxnj9DWAJVC3XyjTrlexd2z5aX3PDWzC9GGGd25CW0jLjuNZ
2WUopOCt3lXMUsUpKhBFn/lp7YgbjSgsuapLJ9wU3uCWM/iocukTxtVnRlJTvPCT
5Uuv534Ue2pXijgs9HKCj6LZko3MGjyNyljUTHSENMWGelFJyHzKKK65f1NXr5BG
hjrn9P1qaR2yWmMndQRy3pXmAYMhZ5dEDVyicQWttoRVEGt8q3jJ2B2DNEpmslc1
t/SCH1NQO+K5pfQmR/O6bTSTlz/TsvKWQuxr0r1EXHGUXKGN65leIuf91dTClktF
8BRwkoqPbGoD7jca7GcpSGEwMsrZW//gmuGzGStr7giuW82eySe/EvPnaKnQkpmx
//glDPZWhCGoF+NAuS/lGWsVImj58zADdFY6WP1zv4buBSOfp59zZwp5LuvJzFjl
OezpaUf6nz3wmRLEGI8XOveGUun7lEN+9fGP0PacEJ8x8FoiP9wNxJUj/jcmVNi5
qTFSqZYQApUx0l4+6r5IRrTmXH01KpHkhQyzB8AVOaaRgyqqMmOD+P9HjcOPnu5M
91X6/LbK+Z2MIG1m3vyeI+zX4QTCer8vN7+wTU4azQQjksCyUMa9hTkFCFs2w+FV
qG3yL86yW+HHijs2WKn8z+UosjJgxh65VCBkO1RpLhJiH19qxOr2qRW0zmYyEEte
11IiZYuKNMA6rWWH9TUfEDQWNnnvIGuTM6aWncGyKns7ElKDlzpAYDBqPGS+aM9w
peyfHaApHEUWovb6jKfwH19PlDSfVIqkz2GrMbbuM/TKV2pv7svcUzaF+FPLHACb
Ql+5Ed1IuJLP8H9zqllfC7kyNid4ZWpU9gHILarhNvhCAQz2xjaKyJ5ibwcHRLBg
LW+Jjkbw3ZEkJdjRNQPa4vIafiF7fGebIFtUK+9MhYk6zPkvHugTPpeqjbqsTFag
J1NKwYT81CNNS1f2rVCvFhxzE+h+EZy2eKiuGj5PYngyQNNWk8EV1UuKF9vx3Mfe
bZK0+/SvunjCfxR4uWrXz4iQh1m0PLZZHyiL7th0uJFxvVBRbs9YG5++DHzYG9tg
Y1qRo3ww/ANddmXBZKAt3EH8XP5PF82U4HghuoexOyxEUQMw93Zqm2QKyuvhH7yG
4TLllDKOKHwSLU6ROQhtsNXUDw8alY3pgC8JKzAEZsaREVMcIULCJT+SeVT7Vlpy
YdjBDjmJfAdVjRyUFjK76954wLBZwk9gCgEmH9X1MhDEprxc9hOVKncPb1cwtuEH
AWEApzsGEc1q+C7jIT0Pd+T5a5Ddk4GHzP5rJaSYbgl6dC09wbpLqEimyHDINaAg
F52d97eg9kSrYsDghPxHtkzNbmmx6v8mdnMGkKiT5MOO6od50pTwalkVjVQwDtoe
sI/mMQ2fQ9TfvsUbef/YxEJxzQjXr+OKhR8KRHHsLm3LN08TTitjsM+2fZpkPt1x
FWlYvlwNcWun3e85qOeAoYi9AWvm015HrxEr6krtVBELZrHMAp5JzZKItSY94wvW
3OoaDtDhqEP5o126dZ6NgJzNLUV/wSPI7hjLr6O3rVd27K9MHCKHwjaHl8hImp6Y
0+SOd+JyG9d+NkOIoHh6vAkxhHx3OfZJIEq/G8cYgIkI9ZOuS3WKMcSf1xBekJt6
fDgy3+gih9LFvOjgH2TsGbKvS1GdLGC4Qiv/T1kO8rc4c/t+xfa/KJVvwEEJbtRx
3z8C7tbWUk84f+t3b645Kd8HwTW/DmFOFQXkzOqFOwsO9FoAijcLZXnTBgKbA2m9
B84g+GZ0cmKo3z5r3js0I3nnK0FO48nz+6nTZMixo7SqDgurNnuC+0y5j2mLywWS
lI+TV8opaXRE4tO6s5iFmlcHe3WcmRJrstoUWcDm+CmxGmH67Dc8uvVRy9l94NNb
j6zsf66arX/H5YoCiHMchAOPF9qmPb9bo2uJcqwL4bHgpK6oldpMxMEYgqxlcyRk
I8LjWfsphtgi2c0vEayiX2OJXd+1qy+YUlHR1hAJa7OHDHNjctSZLRtnuFKs8CyY
oTYCaTz3rd+O4VIi+1CcIZ6qmWcJPkBh1+Bm9cCnNAIzvrMrlM/fYzzMMyEc3HX5
nv1YiZgaE0sBOu7SmaJX9opVWm6uLhiM4wNbe5/+0NOr80VgtQAA50d+wJV4nMaN
qHdHC5/rcLMixflaRo8deWpdhEMj3M5bnkqGEI4ihn9gpKkUIg6cxx1ApMMLk9SP
IzAl9Veuc9DGVgIJ/0a8Rc2u9b2tSKq5oxcLpUA35Ckz32wBkoWkVhlJ3v/humfR
kJtVc4oxKNIK2qHD+bMDjFxz6V0ZXnKcc+2pa9Bhsbd7vqJSUejnxisBc9XZTieH
z9tJIKXYp7kwKSUdE5U7bDcVtw8eypLBEOWQRQnO4CsmBikAxKCpjA/3iLa6+LUP
a4el/6fvfOcIVbFMepac14wp5OqitOZpy5Qk9NSYHMs0tuorrgeZtwMnL1qTUbMY
CRYZzwmQXClrOB/2TTGK7DTAJj4gxmyQSG5tdC0TWsSuP1x+/OAFImY6vMb26xrs
x5n7t7b+CJNdUc0NUfF8S575zlM2p6rYDSXNL/WCFG3dCAN5DxI4TNHhK7YVGkrc
ccQMArDzMWjwnVERHGTgFtDjnyDAdAXcozWPJlW9HxsCL0BTpWPdcEbNgnDGHO80
mVVg2Nvg5n/Mj5D9I6GxKiLs+8RE86lgsUrrm9ubwp/aMsfcJQ6mT3N5meepuf8i
y10GkLKjNDLGAHEi2uNMyisegHMXh7d6ai5kIcRNI3j3rdRrIdt7JsNvZ8BScGIa
/2sOKlChnVRUgIqspaovFc0fORKMISkwbHxLXyfWAi9SKjTHGGsNf20sCAidVkIU
qzQ4TqyaQR2tQ3SUohc8GCJm9MI/074MxzbTC/Ef7frHRZOzVSzWZRa4UqUQOLce
+FqYVGiN1ONGyB13IftukFHO9dpN3JBk4089zG1ipdDzjKjizHaDP9BWHsca1fzd
KAuG6/W6AT9wIdsf59Cf6hrqN1W1Nq7OufxheqZ1FzqcLWhGqX6ufXrscbnLmXmF
venGYoDPyflO4Yy8gj8TK+CW3Ck179ZPDBPK87x/nbaDVBOks7TdQmh5NftlzTqv
Vg6x8JbsEc7mQ4Fvf//6U+u2UUhjBdpSYxX1d5pCHiZRWQSs09WyRJqOnBTKbgM/
uyjHi9+fAX0q+bQg7dBxP2VvdAMRlkuvR7E9DPA5MhaNLOqak8sa5sM1aycPH3wA
2OJQxWksnv2cAO3d1dnUHLuN5odCH3TOR8jhQP9L7VeISW5nDU7bOjL79LpmHvQL
mADeEkDNjVSUHO4hesofnd4Ef1s7rwGYhkUMVRoe/hEwaTBnyunHyUnwV1fxGWnX
AlWuIrwJN4KY9dRWiddfbZ8rKVHH4tWtQuq1VWAK5A2b/E5gjIK4g/EOPwBI6xqJ
mCserYpI7ci0gra8/bqnyAQSesMeFwUm5QdyoNwkRNvPKsbkTqn3/pHyjxtZFo9n
zRTbLrjNVotBlZpunJGY9n9q6vvyiQf4P1G2hPwRUCcJgq5gSCOKZmFAqWraLSSf
58guUiVTLHGiYFP1HpH7XDYHKmkgvCUajK3TKbjunLEvWpZtcWvInSzOMwTujZro
FZRl9dErz9z367+0i4w9gGvRS1CAzQLmPzfNZDJCCDus4I7yN7W3RlAvYiHsyh/E
KlEKVJfGTDTmzx3jWZy56IGaJj2A9ldeOXeBsUhjmqFSTVBLISURuzvfGS1EQYZQ
ViaYTy1NN9pnpG0v+NWxaeRFcvL7hoGr+wXDPXjVGfEBg8//sx9vYvztS5XkfOWV
qy1S86Wyg1ZWZrL4p6JdMbvuokG9POVzbGDXFzWjgwy/uX0RsCjVobYpeSKaDzLA
4DYlKhlNDkIkX5SrmGT4fC7EXVITl888KL2nnTHRCen656E7S6yCEjLBX1ogp40K
D1ep5SbYYaCB1tVEObF3WTICovFCrxryju8YxqN/XFLtgenuNTISyTUBUeFCQGOz
he/q/t1qF0cLPOAdGPuxgDE7pt063st77bzl6qV0xKs2DvoDGFLiMtE0bMLV2GsH
BVBPFi77rrsNxZmK+AZCVzrjibtl3LCQX+yLIrQdKMowsyaKJsgGqvxYlPmfnxOM
64Lef1Wp1RK2/HflBhgLw0EiE8Z0Tj6pJqVrlCBOFHdo1wwmVGnKBTIt/S3mKFUV
pwJfsXZlFG50VCYiGTNCKDFMf/APFzwnZK82kmDQcGNrQOyKh88DIsZMCW0GaINM
3Z6UjqSgoqFhTtk5PElwWVSq1xYsteYA1JqZ16A6OyWeiFXnnt1qXk9djGjaSO9B
Vt0W4jqfclz0eT5rKaYmg9gs9zJerwBQgvq4VntWQp3cAtgu4qxuavdrdt7lr7rD
GIscS+bajFpKyR6usGuArmks0TwVpLwLnaS/7NKpnGSC5Ty2rEy2xA2E51e2q9op
Qq5kzxgmV69UwhsghlyIhPVeZAJJfi7YY78mUgIVwzB0kfc+MiSSdoB0HEnDpfxf
WzFk3J19Gl/XHhrmJFajQZ170Mk1dgKn6xL2I9QMLIbbRETA12OeFnd2H7GIqiRP
eRPZc+EzswJMiXNW+/caI8yTRTvhM90SBjclF/lzZDsf1Db7vRgigGal71fOyHf7
5fvAetz/2uUc8KJ/DE7mLATf8c0125+955Tz39cVeEGxM4abEK+gyVws2X8VbtN/
fbIY2YcYFiZCbn/VCdnxLao6c8Z10zT8Z8zPTQL0GyVib9gy/za5gE4EqfB1JIKx
Ox+/mxtC6Ptyw4l81GeTO7qSaQsJEdxcOKgGIAKvIX+o6w3AC0cSS9hUmczcZFRo
95DDYXX2pjitXSBgwSmWrTFaCsvCKyFszno+uaXv9BuK9q2RD+OfdH5YEGU+KjHa
NDNHQVH7lqimcUXdPN1UTfDskOsxUVWzO07ebkBNJI/18WRPjV9hidsau2dtI3MB
sifrBuUcI9ETUGqsqFG8EpVUyylbOUGw4rwoKsBuM9ZBo2WCBXyDUxk7FegT8XcA
PX/KywsxqUlNf5yBIId/wPAD4A8k8T8UzePQxNGzw7CYyKqBmPj4ttNy4YOF8/sL
4IpaCk9jXRErMMUb09ZuM4tm6wQcBFN1+YMWPgfqQDdv2ohFYcuf21PWcM22icPH
IOhlQd5zcScDb93YQIYsnWUweakGyfN6+3eoywJuuYu0nRGjZxN85p+PUiypPT39
uerfvdShTVlzpRnwQ5+z6WhU6VEHP2iLJY4K1UYM2e4fO1REgZ21vdVr0/Y+e9JP
6+2d2e1x3M2Cwd33AfcrKWGyUdmo27kfQvzMWWDjo7cgv40PydQcuHAY44lp+krU
sADPvJ2BlABoyxsiSee3cs6B14yzYaO4Oa8x8ueah/Jyyo/wOGGJog5rCzobjTjr
nKhYcH0ep0wmGb2zkVOnVvQkEkBKRyMXvV0Oe0eXzzIRKHSaGPXy0BKCdjuAuAgD
/dtAQ4ytmATIkD5Rf1uf1EkIF8wY2+WtPdUn7Bi1IWNk14aRk3d+AsVnVHeeZNDN
DgsHI3hL8bj3JxXPmflOaKW6fYzg3/GKhHc8s771Meqp0DMlPpmoxDkVDJoFoVlB
dX4OUkzWR5NdYwLYXmo3Sn791bgR3XOg76tc1LjYjN/y/cYql4Nl2fadmSI2lLFV
WGFTM68pfXwx5SjnveVB0T73+Cd6R3GgQcGP037tsPy4zsZMIwfORaDCNDmMWht+
MOpSYH0fCrUCNteii1WK/8NUQnaBO0zrOidAsu77RmbXYoU0vmPr+dcMjaf8N4z0
ALPIzC33mXBm05w/n3W9ELYO73jTgf/vPVRS88M7+RV4UI6wRwN+8+xoqpIbhMhV
6LjB9QpgUo8zPUlPGNUyg1QZWr4MiZ9BITUa4Jrsaaf6IMrxKBIKQzovPi99CkiN
n6YzrWDQsgnNi4OXuToJvB5YHswbOkIIRpgKBgVZ/jrukn+tkeJQqlkihuTUa+AV
UNuwu0ut9Qsc2HeZdyCC8Gh1dR0iCojKY2PkmknIExkSsMQ8rt32l2vzlhpo5qke
w122aoJK1FSBF2r6ZEiU5KRg3b4hjUWVshueGa7KF8ScUVxrY+bVcfT9saFpejsF
4PSHFBg3FN3iWPtal9gFxj2iVXm0KxUzuO4WFoi2Jp9fBFsRhI0IwO1DBfvN5VZC
+HY5vWJBuw/A8zEkLro79eKgf0QoBnYPxgxdiNAuzTNNtJrXQxl1EhbE7liKdeaS
s0zT+cuNTs1RykI5w+WMV5PN2MvkqagQhssQc8HHxQZ5SH6QDKxLRhazZFVHSbuU
tO7EO2R541Fdg17AnwfUAXKcPdK10yooQvxZVLtxwyrDpD7zNVae5aNfvo/N2GyT
vosckh2K0XD5tloL5kEuTdRo8x/l0wNiCgOt3QvBFJlXkaUgGvwg+zBfeX/grWAo
2Vkk/CZkWh9+67GgbpKOlaEDMTfpcP6ViCFJNTr7zXIZvfeBNOmlAQgGW8uFTdWO
ZjsaJ0uSeE4ZF5kPDcpvbNX/1OGxHRSkznq5K2UTjaXROhk/Mxr6tJdfEs64+ayU
d6RrEjCsUfQHYZIzLpPViwQoObBastcPUPj7aH1Utmrnys0Bw6+b38C51Vknrg1v
D/BoAkqaDffzX+qfD2jyhBszsqhMreEebAKi0iM7D/C39ov8fBYXeUkTn0leJGZS
QX2nITvPP1hHEOK9xMdU8gJ6Kix/MV4ESwNtuWYesjv09Gp5h/DsBoP6h4rCnNl3
x0e1z7xxRmci7Ga3aNBJKP9k4GWbwhvgjoKWiRhCa+/QBKLNtAkn/Y3Pwx0aXQGy
Xx676ekHqJgXpZtWTgE9yLipWWSZMZ1H/720gB3ywL7AELZ593/gLCqWBOW+w4d4
1tAoVD5bU4AACA+hi2NC32YeyOuJxtuvGp6kNG91bYqG+qiVjP1BYmTxjuuK6sz6
w2bTSHqx+6AXJMR6557E5Iy7IhT24iVbTtKYwUEH1l9oKelfWrIajaBtEkKmz8fs
07goCX4tJ+ca7kxjef6LKemwUDVuKsaSjqgj32idefkmSN+mPiKrR8G6Bu2mQoAz
uMyXy2OaeMIa2zj2Wb9v0kWo/Rf1mlz63pINu7qLVFuCebXff2MzYDG9hE/PdIvJ
tqCrU5V2I3YrfuxU35PKKlmTT54KbzYUiMk6Ln+5AIRwirOnpycT1kwSpx6YTZly
JYevOqp62rjzRV8Iax3x0UAyalEDQZgF6RCBwv9b6IZI1y009v5pyrSRgXpRwLYw
XjmPFUZUTyr5yTwKEPDHSfKX7XlHuqSuZ7L0r8FMU5mZdDKkyAL7sWkl5+wiqAka
ynUynCm1p1ZyPYcVPukxM3dGdXVkErdCk0MnaA26XYZ4LQgMoDs4g1JmKRFhq/BN
IVCzUP3HBxDZzCNL+uevQ2TVgOl9TrqYVr9CIzxDuzHIvu19SaBDW9ndNrJVCxax
EwbUho7lJJANQ5GSvmlB4YIcmwAJ1bMiLaFxiOlBWW+ZJrmUixeZBOlIHa21kOCO
pgF0qc39iYLxg7hTryw+Aq91z/Gsd0aSX8uuA5WCYcF2lfq874aHfTOIQL5RtQpe
BtHEMRUXAiwnhs09TX7ssfE6lKRw0M4JJfkd6ONZBuCms7o5/eehwjajV6xYZ16v
9Y/DOr1JzdDmYQKcYBq1Zo2AyZBocaV5F9Ww/uhsHwB3ESn+J7QFkE32XxvOsiWx
yHTU7pJk03hryTwOJWdUkqQTsfEYk7zs9xNP2pRylGvwZRovuR8qRvLSUuVVZGfj
I8IxYjUwMfsPGCCXIXb9iCsLYUpv3SqQemKFpCsp/K0+Tm5Fx8+6XWoHRkn/6owA
rXMnW5zJZlW/OYgSjkc9DVPXWH/WBcBPh+QXxBoLXF0ixXfu1bT3wfRSBc15vive
Bf56BxRhXQfN6EP7JFG0umLD5DcyaMmUJAYFcgA9x3qR9vQqKX37YOx9Fii3jOZa
fTdgz6laWwqfV+/Io3t8heAnjBrvRBvPpr5e4OnsvMrraqsP3pYqUgGpVQV76Q2K
vWmhyM0JlC8XMiCmO/6wtiz44XToQeIK1WcsG1DvzhHRASjyiSH/gKIHBCNWElXm
eOBlBuZuA+/qCbMOGtKu1KKvcySU8r9wa1wzO/K7IzBrSZeWXU+awqQZUaDqioXb
OALdWsLFwzCjNrSowfhCu7hAlYCK7/dSn7rMXx7GjnG9sZkCViuEF2P6fyTMujkW
3MHlHzSuzRFF5gywS9z0X1cejU8uEldQWyWCt3a463losqHyfJD9vmDuBY3coPe5
ClKpfIkGPoyOVOarRKVzp+zGLjHExdGChwPTLmGtOUvWqngfK1vCLAT1n2ovN52D
yAbNo1fxESMG1ovXTffR+IJlEc+kBXJzxKJx2j4JinotIhO+Tqai2gT3NwT6X/9q
cPmm7r0puCTHMBOj8whJLdvDoo8cGY/YpipBLQ8ArxBSi367rGWhTTqWaKJt9oyQ
du8Vm+x4Gv+SIdrk0r4WJ/Uup7wrDy6DZtfOo1AbCbW6ghCU/C+zTPJtnZPZ+fIK
Bw7BTznJ46qCVMeOZIQXciZsnDdDRtRXBGtUnQp2Hv9RFahdpz/qluIGXjSlR62h
2Mymo/jIx//LtKoTXRaEPsz8lXSBh8LwrMh0Z0h9G1xuSSrnzjRYMqowmI+lpmvG
ATAjxiqGXPNVw8yalgn2NNGfcVCwkN24H/cC5BO8OgipDR8Ya31IvtyJuMQwXsBk
j20BVpDcRgquYygOO/Qv0ZWgJi3TSXJrGPi4JQlfLKaoZ+iIOlYTTfpX/Zj1Dg4x
0wzipniwkGHFZfq4QUvYBssziHI7xQvkT8osy5AKR1X8x8RapyBtxFEBWkKa8+FD
ULUnLKf/U/IdCGqOJd3EVjGp7GJxo4ApUIh5XhZADXrUSCfQUdVNJclzBRXGrR8+
cFgeclhipKcXcW357gZDLdpFh9mANUmIq25ykhvbXmWN6wjTywx5JgdW8NBNhsJJ
VBhSgSAdwuvfsJMwg6TLf94sZc7qei7Kk94VcVLm7ykHP4CVxS9exqLuiwIAD0qv
btUV+RsBV2jbdfsuLYd45yONAxv+2hWXFFVIjR35mjdeumCHbshGu9lgALiJfeCa
FH74JzS9thNa8ChbXTWiLk3lhzoYwaDs9frJS+V9taqpX5NpQfCJzRP7QZHyJNM6
wXSs1D0G011X1CRggqzKOcg9yHg3+uFF3Fb9SV4Fzf95qFA5ehQUVwpfw6oRAbbF
kqN5pCIWGlhuDHX61Nt+4mfCbzQCJHt6euXaFxZS8j244yr7kdUiKNl9oUJBLGPt
KjETo5ZFc1aFfFVmIyupD1TM84NDpxuc5Jl6+EpamWS5ZsrTLaxKfjRucfFhx+0j
a+3CSP8dNylztUU6/BwJBrRZKtr96BRbd1DhaX1MWOdeibeHmReG9gVv6FI4QqO2
zpi4X/zCOTU873M2RE/7pLC/5QxoH93vCsCI1FRRgKRKLUe3F3aZifXVEAtHUT4L
iLhZPRw1uiaQY9CBawqzsaU4icp7AuloBQpGMR8k2NZtkIEkjq9S8sZvFqrf8LFr
4gxZdINKPKMe9D9X2XfLvTcyNjQMXIdwEp93R4dZVLpV4j+KotADW5riMxW7RYWj
Wne9BW+icRBeOBceV+oXvDg4Wu4PGEbdec7F7PyqExVTqeVysDe61/I1etcjTTJb
wCnpXOb1sFLoqN/qnxUOxq65XwWe2SFRcUb00tQ4aJwXqtqyjGPAAkOiUIhqjdA0
eZ5cKC7+IZwp4lddbkl4BrOEHrq0CWRTufE4DVI/l6Oc/SyTWiYJaZ2tWjUigHD9
67aiv7qfUAF8jxYr7ZCzhpoo5ALGKRFCfC7h5YtZT4Cph7dyNtecWBybP5cBaq72
CDwV/4yhcbkGsfWStMSMLt6TRvV1Tbc76zIChzxhkzp6AY4Z/OBYG6qlXHT4f6Uc
RcCE72+m9XIluKSPDKf5hwOGr5bVxzd6thVx2C+0BdK7M87niPvidEYAeR1aBEyA
Ags8kVF8D2ZEsBlQE7ATho4MB4CXtNiLRzonuYoOaU58Ko3h96wSpbl6v9VTIT6v
y8UESH8WvGSmCsyZniBcLISWvnBNLLKh86cTgCYJv7SF2J8r6Qg/5bJSOb0TP4pB
OWFTQAAGDjn5TXB+gKfZwlY685dnT0GlCiPS/538r6KQfA6e3mXEe+Fyj5dqbaFL
w0lxe0k3qI5/y6BnI1IN6mUeHqLXSyzGfwYaSIdgem20xO1qlvS4Y5uebDLnpnYr
3rkytd5+lIJuuuliuPcIVXc4k2jo7lRmEjUmEXjX3PAFNWhIb8kE/VBCThIOY5yb
Pq0mi5t0a+h0rQSzYczIji0eSLXYB4IgMTU8jRl/6fOkEYHea8jcganiKfgcbM0w
4Ccr5MKAQQtAc8ui83ENg52lAR+wS3OflqPuo+W1AhCzChdjPdkDjsNy5Gw7r1wl
kxirLu9bUc8UFISaLpSX7fIG6IiSJvYMXhvLtd1sHAI=
`pragma protect end_protected
