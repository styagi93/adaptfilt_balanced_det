// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XMKCXVvaSNRWK7AF3isPdyIjV69A3VTGW8PpD6RNOUXSOotj0mo+aaqmboe2gHfI
AQhWJZi5oLuv6fTPrlP6JVUXnXcuCCym0QDEsk2Nh3iqRkBXMSxRiP7/H3+Dcfbo
wMBppWQ61MF3Qz8adV2PWElQwCa0UJCPblRlyWD0Psw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21312)
+j/wshg07OTDc4YoZ+9RhlVLKhPpNj616zsLBCN9Nr1Fh0rreLRtni+s621tZilR
pGh5PYytO4/an7s5FftOBEMrf7qhJqzi32/ij4b+7s0oPKynxaJeiFjaluvYH4D7
gQKB+VRYaCdNmbcbZFYjgq5sFcdNWm1L41tAIWWFwy/TrbA/H9OJKG5zFVyh9Mp4
AAwvOp6fV83gZSfhgiVEC46ZVdnl7BqoUAIuJn16yZMX8Yr4pRQFRW2klA2jCsUP
wbvvG91flisiNLyJDLEy1WZvvdGDX3IfWkwOgFv3CiEavPXX1i1U564YccZACJrf
eKzlQE5cNUk8P9/BV8qUXcK8Xx4iQ+wUb4ioNI5aAd07YPhzWVuoWjcRn14JUFql
ybiOqwaTVjPcoQXBabqjdaOifyOPK57+IT8671TuXJknGUqNl30i7TZ2T7UpcEOG
F4p0uMkyt5JQlsI+6Tga97pAyxBqmfYmwtsR9K3so/c8iMLFB75oR+8h1Sulnpch
NmEDuWUxmP9CCP+JXlsWdgAm8yI79rH9UNv5cq72wIYy/eDb4SbYWC1qa854V9RQ
5ncjpI4N2BMMEVzWOtJ/OVSR0gwxLU2Q3bVZ8LSDcsxDFO35ZYsraX8R3n8TG3Ku
K3i3qUCJ8g84j+xgYhKamUb5tUNHm6/I0eBs1ViusYpXXqMmOEAPDKASWLzIvHrd
RAYgQISL9JFgBIDUymV0GmUPa2BK0Cptku8Du4fDkUE6Uzhz5nUi7msSc0S4ZrEk
T7eZpYxYznaW1tsKXeFVeuQnaiIqipyfJVEniQlPrzMYHTS5giy7NSW/sMt6QVip
ebYWNVlKpBcfLffACswF4aPUYpb9UHD8JoykhkbT7L/yXz1ssVclvYaRY60JuoR9
EK2bcBD+lEsWmQHgI+RSfj+RUzx1gQopDMOYZqKwvXpZZWENdrlJfmzgblR4ddbj
tWP0qr6MttXrKk21uOcPBnH66MJMrejUzMIOx3tChRreYH+NlsyoG+rsSb9z0VD5
N0bjGOSEJh9DviQBIUbiylxpTyDFV8G2pNbJPoD6VbS+dZMpMwV+1kYQEdMcs9o9
vOmKa/mApBPR/w7mXz84ein+LDTlGWSI658VLiSXzGjw5kGmGBv8fneLeRCB99O3
7W0TUNQOodgOwvRCYeTYLcU3HD+FsFtYYTfh8x5mAfnUZE+jlxX/+XOnRWRJomzY
ovXB9YE3V1e2c3Zb7i2PFYdcydxsQsaHBIh7e2CouKjPEEv7KMv5iAtBstHa/MfX
KCESoD7XQI9M5B0PrDKYucI0EtGboGP7HwtFQynh19mtFM+85dc2Ye3ZXgGMDiPf
2rgnGEK3eeKnOCNUk0UUCWbUlQskHxRS6JscNyFOQsAGAtU6SzXpqE2LiQ+NTuT/
YKvAhA46rZl5m0KfhfbkBWmXOXbvShKvdPmQKNwwNjTdoTlUwsvxkrNNcuFo+Xev
pcWOh/Ic5ql+M7/Ydfo6NPFncguND8Pmm/M7/CtI4xacdQvoqqP+dfyCKZtr+b6y
jC7T62OskmB+rME7I+94HWBT6F1c5zcolUaNUnqST5WfuKQojhLhCi2aruMU1E6W
V0KkiCYHxcB5Qez6U+LOMGdnOLOJOKGTZ5go5oRXwZNAWxjTbGp+NTT5arU1Ao3y
0qsBbKdzOP++vmNVizTTVWtOWmfXjViiAZrANTuTVfFfkxq3aAI+PNS4biLTRjsz
RgWYj4woYOj5RtuDdjOn+ovUqL2LN00BWcSyK6NhHxwjeWy0aOi4xsZVD4g3IvpX
zvbqThR7ZDzduKdlXxzWMLPYgxuFU2PKc2mkNJX5EEuHg/rjVh5BdLX6n/qVwLQ3
dw7I+TR9CSOGI8bqM6YmtqkwP7jEWKuNVk+lfWXNVyejlEIqK1D58EEJCMsrh+TX
2HvPKqZe55nNIqPIY2r1Po75Lb7lbz28EHIDnJ8SyUqobKPlwY1uzLVsitfpTWNA
MJ8NJhORMiIfo/s8eVyLNFngj+vvosc5J9qAUI97JXcBBtPQpVjESTgy0+Ozi6xU
Z5ANXs0edHGtyc4XRyECr8tBf3j8OoZTPUVpxL5tACKZbTim1yIi6eRpiBAVa7yj
W9/lo06bkz1FVs5hLVRyl2WPAQ9YVOLNSkGNhwfDVo1QuP+r6zSgqYqwWts3f1iw
qEFEX04Z5TUlHMBuzOG0g3z+ROh4CW9mT0/E8biXJgAlz4sxoq4npGJFnOEQth75
wFR2b4YirumAX1zxYAU4TRRKIKZbjPimYxIkR6b9uXYGHlML+P4HPm9gtIPozG2H
oTM8RUdQ5hXnZ8LbmMGKXrh61Zvp/c9PcoJKjeDJnhd6aYoLn4xp86ql2iyKECBY
He8ED0aAi9AdrFCZb7l/baNmnS3eW6HMafE6IdK/ElTAu+x5MtqBRlUjLnkcSWit
SCPo4Dhp/y6QAiXwz4ZeRjVJKpLLcCKhrpSm2p0AzP58KK5uCvbLH1rI2w8zo0PF
Hbjy++oIJtYOUfHjqCWSEVTtGAwAkuOCQPyxUitcYScevnP6uNRqLgPQBPylTROB
BFad4G+ZQm3WQpqGjEe8bPBy0dsDwulihDTaQrfrH5zJswM9tW+TNBrMr8FrmBo6
jQI+0cWS4m2HdSHqK3QzwMDNktcTWU/SUTQWozz8/4ZRL38jTLpMpozRn4+jDmyv
Hj11mcyBnRKMMk++JIy7T/1YWxMW1hsrJhHRhJykDrrWigoqQVQS5zbhUpeybC7R
feYonO6WSMUIr7gVlJfsMPYKNSt/H2qp5f2x7Qhmmv4zEGpChPh9jI/tgp9mCIn4
vsAc8rFI4wTifm9lczt04bgVKCkMFczJ71Z9MyDKOmypRfo5d/Jm3A3+1pu+o2YP
mN1rwTT9TRZ5d/1aLjzRQoe3hBG25gVSQWO6sToV6ySqcKk+lnKUOUF/RgVXQTou
5mna7dfNr4eRSSYj1aiB9AVjJ981nRfQCHFwqQW1gjBJLoPFDYfcEQMkTO+e/85L
VbnMD7b/t5z+dUQK2yq7iEoGEiJCIN47zKScaxAP6FtEFmr53Z6UAFhWbzZtBlgt
FhoA9DNsyrYvQalpPw9K1jKM9+LZadweMSQCET263cVvZLESY3Tx8I98Ktk6Q3s5
FQF5Or4I2TJ1vaScee9XkmxUSGltAny/NGnvPCXYuUD2q/jdTUuUkh0eMAdhmTJu
SWfy2vK+QntePvKacKxM/5n/z8mVdKhylBWEmd7NfZD3b5yqQH11nvB5ntFl73C8
mnRGBgnMkgJyFdG1dJv7n8N+mltvASr+UbjMgno6zKXqmjv234xa1EKnWp8sFctp
wNkCcRTs6ScF8whRNYX/xS7OSPeigMqggavjEmwqpX7Kxt4bZtn97YycbdK8OeUj
i03nJE1HAm9NmiMjt2ueBBzB+QaDrbl1KJhFKkFYYgkTQIxdqA1LPCHrKIX+cSqe
DZ0/kNjtoadmAg7D7CzTxr+W1ZT1VU2YfBFz4o+kpt70s9iuM+rX8jGBs4a0kpAC
9ESXqcCKsUKFl2FCNTuiEhCZU7GIffTom8UHVjk3H3oBnPcI74Wz03QUrxTqIct2
06NMnw5tpl2mhQjLKJ6gF5MfWcww53MD74cyRAzfKrqJaAGd7vaCzh7rTSxbtBsN
rd2bLEnjV9V5b3htZ8bhRkA8aPZxRksUGbSEIQkpxGUs6rHeGdK/H/cWA/hhrNDT
vlgk8tBo3cwo3Vx6qqQyCwQazooyHxy2vk+aJdIcnElgvUs7vEvXS5EEAgA2+aYh
pty69xb3LAkZWPmluKzwdJJvaDFWkKl17vhbxmk0ScvHXy8D5qsV7IKBSxdu5aK4
QWsMPGoAhqdfSzbzYd2XpbCrmVq3vjx8AUe1smOqCfJBXJhPxb6Czc+WSMpNo9dn
5XAdziNTkW+7uyWBL7YOk1kzcGECB/sdrHG+lf7zySUdjLLC2HKn2Un4FpwHjr2V
nM0+vE1dFLNPCde6Ylf/pLdmnqxV7hn7cUQYe+9oU/sQeDv5jXFQO0sVGZ7ZsQUZ
25Gbpba615p+iTiHF9+wWUDI4UOQHFmidMWowraz2XDyOZVutuQUXTB5GLfiX++I
TGMEroeUeA/AHUipht2A8lNkRLG3hE6+tjlsWEJ4QpYueD91LUMTbYJWhaC9lL55
9B8tOecZBUeNVIe4D9o3jRsMy2e4zEsWc2hTDx76pl1FxLY9uJik9Hpg7kmsD5MR
Q4eIVCJ6Ib9m+v3xBwoUia0M5oeR7UqmFL2mgeJFKkZJm52R2AWdouumjsYl8V+0
JKBRCiVxhaED8gyToGV+caAfVrCF9zACwF46oyh7/Gf0QO1hG/fIT9LCbdd0vEhp
2iBzulq3QgE8GdRrgwwOIyl+97vcKKfdsFrNOXgTe6yogr6G3yuV3wp1s8n1saAz
KT+XsaPOxruLCVH2u17ERvCT1sOjFiV/mJIQYPkI+ExcUGCAfiNBG/oPTAVnk5yF
q2FreQnqIV90FmFYZnSsDMoguGIfk9HOXeE1m/3hVGegIfMrIN13My+x95nObxob
hOagWWNnhYE3owQ7K3SUmcvnwMArFslyw0ecL2kq+fXPhPCJIypqUGruwhgYnxVR
wlC5QJCf+LSMVuH4usd+Lat71q1kIHFSvMUJh3iNxbVEgO+wooVqYuoY8cg8Eki7
9kLeIiEYPT88ZXRoMs4/98zJV73Cw/7Oy4o6MHliZQjUwcS7d+Hyt23plj+CXcQY
q0PoK2efxmJBzm/lC0mD6GFW7236KeBZJIGvLodk41Kn2zFm9ycINrwD/zeeWmwZ
cuq2iy+R8gMkKCOgcJgw4A/mm0PAwr7xsZ5e28I8qhcXOyMO5LccfkKGFe7AXXaF
Ma3UHHg3Df2EPsEqyat+5aTIU+33SYDO/bxPX1u4nsNBW5RJJeXRtCtuQdahn+X1
zdfVY7BfhU4FL6wiwT5wv0i2qAYPxT4ZO0d6WrFKz9oGwWLOb/RQpn7NSdYmRUcW
4Dj9kFhZ5CdY3B7Q9vISkG+exOv2rc90kKwKkCCWRnHJDlDDFoVEi5UjI/kF/R3s
4+FSARFO+RkDtuEC5mogOaB4eglZZduqhcxgs8PnXfuV8IbviLVHVNrCoqNWlhdX
HFmzgjrGiiLMB/9NnOByS5G780wvgCezTabNc9L5kcsvrDi10bCG9NHitAUC6Dtj
vjPC0+gFaGie4nJ2eQcBlNMQ7bTsKi7gAwGD/+26qcGTBFipcewq4IrGrIa2hFxv
NX9CRAwRKC7w7y8W7xFF2pJvZTzCrHFu+Wyd0atKGYyICB572Y+S0jKvjOa/d+Zr
AP+/31KXQOBGUs3ziADElJNDHXNGkuz2R4VGwLd002Iq7NnOUpG0oBD5/APN19PB
/liYb/VjvHjfsjiWVQlDm4G/8B3rLMLgYMJmpVbRgzAKkGouupKTgSWtHEl0ucKa
7bbuUsxxn9F4KU/DsWHpod0NWSDvL5Oe9NifBGHNFDUj171ZBN76zu1wlYCq6IUf
BNfZkCbp1BfcmJqTjAH/SNBIoDojEdSCSgJY6smyQvzbBqo/jC4WiDjDsvR/G0ki
+MIpQq40Cz9re8vH3yvoCj+VQYeIV9ypStakL64zpcbV3DPDBtZG2ixgVEsjOWWy
1eO5K6Hu8ysd/2UzkIeabvQ8IFk3b77MWeWbfDA9Ai7XzP5vZdyc0/XQS0qp6e6z
sOfS5gxSSq+Xck5ZqpYAMWtBkDuHkW9xlUJcqEWtmurh8oJ5Kma6YJK2cUQaB7pc
AsARzFQRdIMTK+FUzBpRq0o/kdzEJO5DlAszxWwhVJev8GSH+VP1b77b0pvPIR2B
ywZft79d+wc345MCb5F7mBr/KAylN9DQHBv1aQU9kw/CbtcMFU4IZk8WWe/R3Oj8
cASI5NxvXV2JJQvEaJ4ekI8UehaDoXr+f4dYL7HgFIcaWwjpbzJL9AplQpDz37i6
3vKcI1/obRkFiM05v9mX3BRoOM2DUR2XOCVFjvqzyNfMGrqU3rIwL6PgwvMmE0tt
tVUQVb81bvHWDj1gkUwzU9j/qK1nX8QccsTb9lfBislduI0RGCV8lQ2qURG83u1m
8Kq8ZZWrysIwv+nJs7AUBLj5nMlyP5ie47Y+k46kX19WHD2kfUasawGHtFUjugKU
+2aIdGsJkFJe7Yt4tf2cWkQDXO+uLEz99hf29au5AnexRRyWegPUbLwJvaDuZxZP
PpSusgWQjemSm6BWbRTniE/NpRQ+DAYnD2qnqbuFMibTCM3xj694qlUw3zzzJArU
ZRoMSvTnNwfQheA9LDXG9SuesMhyZk3zLCgClWF1Yb641ZSB1D2b2O1Sw7KRhvaI
Dt0TURmZwT2ikZvBCOgfNytxasMDSRSR4L5ZB+mkRAM14NxM5N/bkA8VFL7GCO1A
kMb+I5RDq5m0S3NL0F3Qy7XA/rxBqf8D/lkUaskyB4pEZYOTAmxgwWqxMcH5BND8
37+jF5sd/c9HYQIRznhAKlBRYeyxUTrAPewhoqr4sTjcG6SWvKh1aTklNNbEvvTo
4GfLJoWCVsgazuISpsybbcm77XR+ytsrzIaMrpKbv2YDtXCphY9+aL0s9K5A53Bm
ZOuhkVDih2Mcsm0f116fxLAJHq7eIQaqaAkMJTs2jnXsfg1p/I3Ww+LR+uzA+DBN
3+wbCtCfSMl1gzrUWmQUod4Qm5ljTuNfmIkLL8Qjn1zjXIO934QSykFpw5rUPE0c
uRIQ/6EFCYFpcm7KMnY/o4kFXyrVLue2Jbmd9BLlybQddjggeO7V+n7dkrtgDFy+
w9XgJ3fP6M5rEDdbsrDZ/85Yt4gYT3XEVS1Sl/F3rrDHThdtmFDQFzSNDF/N4XJ4
ZBH6Yg4FTjuJKUTelKLTDQYu1NbbUR6c4g7Xlvv0EGFRA2yex2uLmXAeaI0HeTAe
jzy4dXnCrl5dqSnfC8fQC/lIYamfaA7y66YPHXego4T5qhfeNiHMv4wtSug+Z3kf
KcyhDiCQoh01GKA03NksLorLgmhhkScW7NJKg4GGcQgpp8fX+sy9qx3SCMUG7mTn
pR2NbXPoqem0EzpdmcyByjCQ1F0YYzygCgnfQOCgon8Fvmb5zRdJBYsraGnLWzw7
W2jf9T3zc5zBkTfwuqbDj93KtUXekEVANU4yOXXPeAm+rGPKTwN/NTNfBcP49kDd
ql/EipZrraRV215v3b8ZR8fXN/e+N6BE8a0PQy0llNPa3wz012xTZ7rnChfFiCdJ
L8TEAPcXipGY9pcmIXwE6kzd99EOqhXk4eI3P4NNMA8i1HATn5u+w41z/NXlsSHy
0Di0Th5kXbBT3Wo0AgHM22b6WdeGMJNH6PM9u06mhH71DMCHzmkg1HYtYL7BqjDr
qArCyCo/VvDpEMEB4QdTre+NxC2x6CNB60FYJHnnIJ3IUKoTsqSAZI/eNkjYzIMX
jV/AZcl6bafBAb6CCu+Ao+qnQuMAZ4B60EkgrL4ZVmzE//wGAsMr5GaXFB+Pa87V
fY9D3voZ39LQUxWyEYkFp93VounrFkD2Ls1GfchuhMopeoGByL4GPPIXVxhiw23S
fzmjW24Gffvx6hSYtFcMh8aZ0m292parOtW6S7v0GjkBdqsbyQoBfj+dL0pOeQHe
iZPOJaqFiPPTF9D+kcFSolT52qWgd5Mj/6YaM9hNDlENCntZg5AavZdexeC/cdNe
5+GQpMse7sISQsDlNTmz+YykM42VeiVFHcE+DrhRmt720O3ifCSeXcq+pXz6P4lS
QiNDMpCBhD5PUXDZ0jKoMI0BeB9pdzWPOnmraw+kogXdbhRIl6XdyzYc5MeHH1p1
Qwx2Q9px7Drqz3mALnCIQXPaBjLRHBU3PcmOWs6jkKNR48VYM/J6AVxfmhKLM5wf
+uQPuQa4JgeJT7be5AK3onTdg3F933JrlN0gYnI/pDzD7EfRjjanCg7cJSuZmWJi
rvYixBi9OmuVlGhCrj7dugnQ9D7E+vjn17fK01zkjI/ZZiRdQ22i7r6Z/vjrUJEM
Xu3GLxhjVI4ua546KhoN3QjTX9+rZcz9KehSAUgdyrg3oVY4F6CqTThVvzI13d9F
YOW7pBiphsbVgxVaCb2QNbBokr3R4Wu4K7p3MivSO4bN5bZ7pA7uujW92+yFckG6
QLCFRqMZRTDP1/OqNOUqW56zkFVPwmhpqFMdlnaqNPtZN0tGGahXTR9UgFqHlRv3
bKasruAXCRnkosLuilGr+Ejx0pbokOCLdgiqRKIMF8upZCbNagoxfgKqjBpSk8QF
ZuRxf9TfUsg6v5u2qmcAWGXf+H4uaH+ay2+PuJCTb28cqR+tek+c33g1gzZpFWNW
XMxCGwJdRDMhwEV+aO2XR4ULV/3FahWsUHKHg4dFhHypL81HV3Ch4frVILeYcNRE
unS32fJOVHGiv3rfoCw2kgsViRHnZwoN0uJDLS9GPBu7wFtThw3DvhHM47td+89S
SqyTDcQUSSuJoBVzT71Lbfi4aiNZIxqICObevYBlrBBw9xj1/fN8kr5Hkb+NWkxq
PUvGfzS5f/3AvW+cxyWq8+C4Iq252jztPEVrUcErEcUvqKpjphyeIv4RxJJqIdhj
RXj1hU5kHlJddenmeGFcCZ63hfHrVrgycm+2FfpKYQJH1DzkIk7UPTbtcGCIM8d9
1sT3NB8ajAHyoAdXypYng/iYwUe+cmcF7TKUx/vTKdNcugr4E+Os6G15BWFnvS+K
f0LnVGjpJkMGYZSv8ee7JrJLIuT5DprYLtMiXtOuZLrCoEFDir1WurIFBkCOEucm
+j6pM5k6voTVdbgkrCbC9ug+4sem6GI9q+bmS3OIFTWOliGUYKmfKfpQzx1oYqAY
NMSKVdXhf/ztF3lg5xaS99M5jt+KThZS8gzkRrnqEz3U5MVwXvVrTiFIdBQUCPOp
4bL2dUtjwXO6gK0wdB6OE/hOOLOQffCrMWzmF9wmcc7hekPXZyThWcPrbeM3cLrz
lo33HU5ZPeeiO+oDosMvwVmZQ/rhxFLK4qUl28ZuZvLP+q/oyqwDk4xZvNnUzjN0
A7K7v0lOXRV3Wp3QuZUk2nkA6bNpVMigSXirxJBExPd+5xTVE/hDlq3kXmQpQIBz
9smlLLI4HIJExH83QkHVyPrDIEVq23Gq9o5zQkxMhafQKz2Co+m4xo5gaQJG4091
ZppwgdCchxDlPaHoisyKi9gR/b21MGOq9F/C4W2sG2AeRryhHZd3TZjpKiZrCeEi
/lA11+lvo3PwMdMo3vZSThbZZCXVpnGcPptfi3x7swRFG+QTafy+5kUW1BVSjzr3
SAT6Dez8dkD3t6/HgM61SLdqS2Lxw/CJWzhGIyI0zKNNHyCxmM7L7eHoGi0TcnG3
NWNNY3CovPhuY9Ct5obXE9ByOtDcPCuf8RvuPhIUdVBhgoZqD+7mPzgUyOIlcKtf
0tC+a4Vj25BgplXoiRDgkARduZik+eUdsPUXygB64wpwPPvOWSgGDPRP/nwd5wHe
VJQoHnvccN2XbkxAGvOkVvMzsuQQvbPVzhjT/IjmMmg/bF1mbw1E5EKMhGEqJzlR
sB0dMie6hL22ogTSMjpXXvWretSmaLxJHbNW4/D1Sp5YFRC9ka0QWvW5eWgaqBMg
7DdFUiGcCrRwdboeMFe8Ppy/hzB46PivshR/SCiJrpGT/KtjLdmivLcR7lJr9QH1
XICb3TF8I3Ngv28X/XLoKJ4l3GJVxXxsxtc5K2GP6aD8zbfE5rqwmU6X1uV1NZd8
+t+9KrWa+0tEFtHZ9rsnduXevoyyiXCOEMq8K7rPWs/e+H7y2FU2vVaezaNd8UXw
bR5vlMV07IWTsuqXl9wC/Dpee3znx2B0kj+ziZJ/sDaCu3QHIwVo77TfDTLK9yLE
BI7aDK/vjoe30ERcTSbZPHnXNb2gJXSKX1rZ/JhccTbf7S5Eu3DlviMb2TNES/EG
gWj6ixR+P7+Iee2ywg7bYu1vn5C0LwvTfFON9XOE+9Ix6wkAg7aUtqOLd45rw2A8
lJvpbNfSKB0GnMmO8uFniUHppKVVktJtbgd2FmPZUS8iAeR6+JoDmOe4cGkAeh1K
v1IhYEvT1i2pBVg49mpmjwv+kUsich3Ky5rEE9Gw7T83bBwZbur+Ni9A+3eh07kY
LwAZi//9EKCxk/JqF/FPM5MMPulkNtqcQQlZPq5fD+qk3pQ+bIS86hfrYdeek+mo
l+snghtULkdgbYL7oiAyPss+9fbOVguqJIIm65miNAR0w207WOlahrZefb6olezE
bsZTk+ZDIkhh+D8RmFAlka4BgBHAh2QtWXZwz7SafAVyox6+re6EeGTRQK0SMXrD
1E/ltLEsxvT0SnJDbOAKGh+D5T22BWIvzwccbe69D9RSwI9WxbfGzqWYqzgSXagG
CV2NqhSLoIisrmyvPPyQBcQ2lE9aVQ9zGYQ2+mSc0hgP+9rw8aRmM3Rpz6ldhN4w
JYTY4OGT7g7EflJjgPj0BGANc4lqNkW61DaGiyG9A033hzAtWWsa8K2R2dt6MV4R
A1XyOcwVQ911wzzGYS4OO9nO9MGeQ4kICqthsuaxmyPCc+sr6SSxAHuHt95es8h4
tsnU8H2Cz5c8o5nv9n3dwy8CYu+5tMIrxNGQj+nfQ7y6Lb2GawlzPE/apmQ4fOof
99pL3oJz4E3e6eW7uBmDzZlUa3qOemDp4GjKS+6RiozJD595REmeCf2EsI1KL8Tt
oB5T1iPUTDJrAqAfH1WrNJNCWZf0Omqj5ugJJFjh5lWKP5lSBEE1qEjfSvWbgLEy
5+JpnrLQoXoUMV5Q/r6EYv97mskT/H5AAaHYPC2V8hIfpN+FdtrDyeEHfFzUyNDs
wdEsyNiMU0+tjblsVOBwPQKhXqesudSBDG/7ZoJ6yrS7MDdZmUVUJAnV//RuGpbN
tIobiBKyYp50DOREO5/Xox4DJQsKgrQHI/VhO0cqcmob1ws/KEbyIKcOWh9PwbMk
hT3MguiPTOcdf90PrzwcW+ygnZ2U+GYN4rdgD99M3Uh4SkBITNaZ8jbflbnzbDhv
3niaIhJhyx4/kNlmDAs5uwlTdv4um5JVl2UPrIBCfWb8rIbJLREnyIZHwAcobfDm
/8GgKdwNVwPGJKXsb35HseXKUZM/gpFuTANrjwZWFU8RfVUfGR7rsRWYEgVPgMF7
Rf//Xg1B6J/bROvjGs2FfrCYNFFIdon5dQzGIYNONdrxshyR3U7BxaTfoilhQEyE
N+PdYhPDKvzi97SKbOHG5YtYU+/ALx3CX3VKSMVthlbuHSDrgez5+K75eztoOIdn
q3XezOHaNDL+0VXojRgn6zXDgDvurcpowIo2yOaZ1fiRtmYTGTtncEVS4EOV/6pW
9QyqwZnd29xkUHwYfp3FWsAwc6tnBqtF0XdNeOe4ESAFfV1bDE7Lo//f/jEKvk0q
LvzLHZMJ9VWN6MLXY+q0eO3Xlo7b+bGIl5e/Ut0efvW0NdpNtntISBzKdbRzZpBS
HztAfpdKC5Bm5rvNedeX/8Fk+yOIe9C5Htf5Ft/8mNzflASA0PqLFYiUArYIZPQk
cSkbT1CUoaZkwxpnKmkGXkFNZ5UdMXrqoSBNuHq9T09ynQq1aVUHwArYF1sYlMxe
agStgBszSNncWP2kf/Bu+7gtGseMyRHamseqwslSFXOci8RS2nq0jB3QH/73Qhwz
a2tP8fBZ229uwJJ0un46d+gPkfCYwvpKs0NJg+aOOISsgmXgLeadc/v6Y9hwOfWM
EN4raCFAes6H9iQxOhovlC0lbdLkxRpMsUG08dgacngjzLKYXMpB9CKDaNjteOy/
OOl/ZOtIAz0orIxuJC0m33xZX/udt2OIGdGrlGuZ+sES/68nHhvJs0a7dFpNgsai
Csd66j5Ym1eH5Pgf9RYlvjxNtlDfwXvShgT7f1+AbgIOFxytK8pLpFv5nP4ogCo1
3y8CdAVzMqXbdTm4fXyZDtTh4FRiJW7SAg6hVF8rD3iGJ9NDD3SORqC+xAKhlYJt
ha3wF57riWQxjyIC4e4+M0bNZ0I07ZLVPYnafiQ35yeUpPSv0LkJ4TbQTBVDsaKl
NAM56wWiKGXn1mXTfGqDH91XOLAYxudw8Nlc0XGz2FQJduGHH175WN5fOJYNcJRK
bJQNyBkkDr/d5/gpXT33ke471bsYqvPsL0zi2ls0hczsr80A2hLMWEpIC1h5XIuL
0okPmVVhJRC4ZKWP1ARbtc7wHwv1+rmj7QRDMDjzQQlr/j7o3m+W0V0lW7kv2jnO
vNJ5BAIBB8UL0TWYMOOQvzhy9u+BKrUz3hAyPCQ5Nxsyjnz+ppxf7b+ud8vMOt2z
vxyleIWs6M3jRn+c9B0O362x8P2z+lSeyvUtpLdykxXmlbIXm1Mfl2q8Q67oEI+7
5oY1NzEK5qY/6myJ0ilvVo+1D2UpEFUMYdzqeG7U2TVzDySbpnMWvLF7fX7JvEqg
tVCclGnaqDeF7eKEUWU8NhN08yL4tDRTa/Rq7DGtdIcwWnFle2t6s5ALw2MztLG6
1Vx5bcgSNCoEPEThpMpcMsudUUpFLUp8Xva6o+Hx+ryDOuEbblgizU33Wb6GirPu
qIosspVmNRh9V99xLIGyCbcR0HKbKFZhOnRMI5o9z+fqBqA4iYyNaAlVYucmiOM8
kCLw2lwbn+OkALbK7utncBEU1BfobpBZl5LzQbt2IeLyNg4vYdWMULTl7j+P8c19
zClmwRze5cd7TcC2jO3Gd2Gw/a9pVcWbFL4Q9pA/MmI0D7YqKSCuoAflNdcc/hOJ
ToyA2D2SXtzdTlmZqc1I3jjRw1AiNxmpco8H2ANAId6GOrpdonqm/VC9+4hia9jC
v106ieVB5VD7YCSAFcf7L55gQAPN1RGspucKRHp5SXch+XlpthDfBvArygHn1n0M
011em0rocGDHaAKgfCkEAHOz4h2/dvjSBP9+5gI2+eE34PplopXT7sz+1RCoz/B5
dA6iYsyzY0SfR0s4gSt2N5ZYd+/SRDDFd39xa4oz4fW5AOYLRG1xC7OX81OfAfdn
b6hNDXnINi5nbJ2lArWvyHTnKnpwYNmINaK5775sz18mNMc0frcwGywbOmuGmN+E
D7XTid5+UkTdJl+pKE0c4WYXZqLEBoMUiYCaSXmv9JpZNc0yXjZjjk0JMqxPhWJC
+Gpx1WnBkgT05yrtkCj8H6CVXnOfc7KW9OhUoNJlyz4lqcbuNC8f+bZ+i8ZaFgN0
P+5pQljCohHssjHdTFkqXgURpkXCouZgLy5g8vbsz/RI/JyHO4+YzHqBpGvwhllp
g7qDQAPXJN8dmsgGinR0/2FoMNqfdTXcN3DtJtSBMvPDd9DigW+/hGTaLk3ey0zU
X4jNCfCNfYjoOVIpz3HlXsAa0gODmGEvuM/rzaQtqWm2hw/8bApLyW0mwHy8sx6L
IPob8aVPEFQOhyOdC90vycP3Z//1S8vNC6ltTLB/DPnUYOLxRvtEubA+9J5L6Kjt
x55T5m0moKv7Y99Wmz1lpBEQW39lj3PuTgNyMhGbNL58zWBl91odal0cX2pcimfN
dVn5JMOTmHIvx2eEpqkTOsWOrl/ObZZyZV8pd9wUb4NLRbNgIFFUA/Z/N5oWDUMK
Chov3+V1sPI97BEA2v1KRfAenPjleGvpctYAXkPDAWXInXVNiexcaLOhChC+ozdd
DCjLpRNVBQhGLlINwAjPMP7+hIrFpxJo9TST6I5MpYOCAqcFejsE6VSO+vWMgmxF
TZQn90pUA1ZItIYw5yRJtXw+Xeaa3Au8IU1lihLgBwnIWO+0J249nvUDCwLY4KiQ
p2GOvFbixyllE+PxT18XKIk2KHn1cR0wOVIBQvow8PmzHRgsVDqAFSdc+OThws9/
swyIOlc3btIMAk3GvH6zPJ31otwE1Gd31eoAB5+5DrthtewOjR6bCXgN3KwnRBVE
r8OmjL36uuqKxMY7MHH57Sr0+DzwNObkeoC+eIbIJc9cO1JMenvYN/KF1Vig22SE
nP0gIRD5/FgyMIBEufY+o+KqUMOFPACvtgLmUjp812jp+rESGn4+UoI5l35OTLt4
Q/v2XYzdYm7pwBxmQxmuRcbB3jLwwtNlb2iIjJlxBwpLGpsSMOI1EVFQX6AsVSQ7
4qcq53OCcekwwDEHx+gC8sIEYPxmmyQzGU4fJt/x3quO7EnZC6UZX2ObHy/RSiHB
aqSQQ0MXR3Ap5tsXqlKSrD9lgl5TUoL0p1By+KPt4BekVsizfonOFSOousOO5oPF
QFyGM28bgrdPYLPOdu5u9pRNzxr4HWYEjAowCimppEJChSf8iNSTKCf8Qk9CZLHa
jd/+y9dKQQ9hG9/bdr18CovFFiovb3pnEsP0vlwRMV+9FZ5O8ipXCIgchxbxrmmH
yFjtyO0TT+n7I5ZXTkwW6bkpG9EZWLYx5LQm56sAWDTvxXvyj88toMlxcmtHTcl2
yJzlODHZWIPFBuvXhEHRsmGuDy5jMNsKkc9CBTX7R1ept5iW5WCdA2tuFs+n8O0X
LdyUc+PDWxEWPKMuHy/GyT0a/CqqPaPlf+sZ/8EGgJAA3z9A5A13c86RHomUASpK
APVfeghQurL035g0WbdNwD3i2rEsThv8J4A8QchwDtAjwpt+iCRO+xuWpoCiN2YO
3m6lLreTiLSW3cK2RCZFUSDSYw4+wgrFNKR7M/yU7AbsdQclN0cl1gI3vQyi/ME5
xXNRcqp5l7oy3gVGgZr4PD3ljtbXZxlQC95TsFUmVuP2vPi6RwML6dCiyG+YrSN+
3Ko5vkgkdUxfBul9Pl0VmHjfMCkrudfY3h0cfctefIv8a4FZlgiq3ln5oEgHcO+E
1DrPuXpp+NtjaSMmNUyZV8etEEnLzxAT1Z8yTLOL5VXZASUkhjbB4sXeKtwATem6
C+o5LnKOQb7Yc3xQ0EL2Uk7/EqhC8/h1Sd7FCnC/mQBZB8RzWOYU5DYdG8RCHVhB
LwntFXs57pRWVDXca4FF5e/kw0n9ZppjKoWmSs1ZHyrUkeU7bnDfRT/ko3huTWYA
w32oiA7a/uvZu/u6mnTxpCuUhG748xfa8fIQoKvluSRYmsIFjQu8Gg8aYQOLqcyc
aadMA8usZtgz8x87CJRDV5N1AKdXipTcc/jeXPplGCHb/VOOV+iB36xGUoRISdW5
TL6S2n8e5x+xZxTEdabsoNnUY7rqwiCz9E7tXr5NFhYpYiXEFlsk5f4nqJNfgJFI
unlf1koQwN21YDCTo5so4h+m0aNUm/69Z2o67oKwFVEV+llZTzWtiDKEChRxQKls
8c/Ef3WyFbH592X4DBXoENBf99bzRiiCboFfzHOFo61sJoNogS9fFpyzEAzRcidb
WfZV6ZSIEV3Rhmhk1lJrTu9/0LYnNaETPhD2svin8wvw/dr99sZEsWqDLdMnjzfQ
gJilgmZwFqOVojN1resDC9Wrd/RE1kmop5BOQ6RX30Ozh9PNrox8mEMaO0objkPI
cAcAbyVyWvgXSd0R3/a2iOs0w7nBDrR8k3KKSvXTMyOE5JaVh8SmtQaxIxyKy1rj
vSgY9MtFpYlS9FovMvv8AqkTc/vNYQpgmfknJF/sn0NV6tyWqnwBHzc7pIcD2GhD
zktxEyw3U4JCgrh5nCV5QJUFQjEZlNWzbxFlY44Xj6pu2hxSLrgYtidlIiqQpalm
UNwZz0z9pmd7quZkjxXbUs9rHjEXIhy2XuHMcNbS2brnEN8aQGlZIb2ibCqlRk+x
vh1F1GnvKJ5ml035znNdxDVWInEIDWlyTZADb6UhmP5gXpids7crxNxd+U/5JMWn
Rz38ZrqptZ8RhSatSjwJVFxtnMIUGl6UReBMn746QMgwXY20+nDTlf4lf6oyArL0
81acHQykPQ6M56JAGYjviOUs2Dun7IeZs1AR7l0klzyqNoP0CxebEMwH0uvaGgAy
3ikw2NgrzdqkLk0hvcJrn3braAazQkd8Dz2eo1afijuYZZGruGbjSQEcBMovGBfs
1b2PDQExfm4uY4nCmdOLFse381t6KLBa34F3+Vkh/aiIzNhdHikCblV+ebPoFj7S
BsVNZjWWpXGJSuqqUBavnFbH82cdoxhsGIFWcKJZS/I8Vak4DYbHUXoEG7xK7dve
+9uQjkJoTquldyY6LXMbth78M8aB3GLEV3oRWPAzTmv8MhWf2wQDVmuvS2canvhH
VH0ZQ5TKsXlezH3/DX9N5B5U+hyRwaemJ9UWA2L6urPP8JyQ7Z6w0ZCCcZFWjiVK
v2jUBHpYr3tTm6sLoIdWOawZckZk25R2EVMK7dGg3A3+NSiSnn+kzziw6o4NgtjD
l8ibHE4BYH/Hpz0O/X1tfGayTaZnH55tV8GPOtYDYtzSvEEW57EzIvmqkNwt4XfJ
RsH4+g632Lng+Iz2R65r8bjmGCfV57UiCavy+XIadvTEQk4QGlEvDFsjmbamrM3b
voFLrYGT/gDIfVdr/efVhk0fjTf6rQZENHHMax37eEhFvC9ZuttY4+0xSgvINj9O
3vAsVLBw8vjvnZPKbz5tnN5Vs21x41P0+yku5xUyk5QF5/vLE4DmuHbR1i92F9cb
X6xJrEzXoXCnMUdvpcXLbTk/XUCSflNrSERa9T0SIMiWVKi59o4w833Qi5J4AA8s
MbZlb4XOO3cc7QVTvBp9AAHQgzDHRWvgAIVFFZHzaKLTVv+v87RaiyGaktEub+kp
pl73Ttp3j9UaAKhyG+RlfF+IEiPlyhKxqA6QiTB/xpNdRk0ORAWpUXYX7fZY4842
0U4turHbmdtLNCO0OBOZBLDwoUVSU2BtamcEapIspYENBL4rHLUfyEyLI4qad1A7
kGeapaqSVRSjYAilqrBqcwnQmY6G1R4vCdEsHhPaHITttJH3yKnF7YX9HXcVpToK
q35802jP3x8GrcxB5CYvAF0GdIfiIB35f0t/M1iLNxngrEAWGyo6+wtLxIH4wABu
pefzezvPWuFgqGo5Qo8Opf/gZYuLRajrHJJkogAnXZmv74J9aKvudEeB7SutRTJ2
bs8tcT7yzXe4MRXNaGXP9VI1wGXxpKIPxjGeHrI10cu01C3Hm7L0/WNkvf/mAVEM
yrm74Rbeif5pv/YdAvl7rBDiDrzyPKR52pTcxOgdgMsOIXF4isGZwWzBuRMKqxhb
ziAvEZx61IvZnboPTK/UjKWjU7q5IUTdywoN+dGFMxgs2M6WdLX2EL9Gqa3QE5rB
/KOnLkCq9cJCyVMY9lAo11MZs9l5ZCZe8toUpwRWUSGKgAcrX6dw+pcTJ0YxuKyW
eshO3GT/JJIWHspkCC3k+NLa3+20A8ciy++yjnzoPgIjg9WwbmFPj3o3WJafSGq9
r4k5n492jd3ffo7q3JgZwGsW/tdhCOrdpoePuG21sjuD5hVgI0ehTjVbxScajGEh
OqJZnT8KAShUpxamNRfnWGhtXAFd1E0c0AgpjiwoNv5xpPVEMEZqh0ImESuu6jTZ
QzHZrq1hp7cHD2eGMXNQyat7IUK648ndZv0prDrrGP4l9+Ud8bRqD51Ij+7JQ4PQ
Y1qKxO1Uyjs0O35m/04Vj+9C3R3UyAtTnhqhTPWtRw5F+bIAnQVpRvWUNhlJqO3r
XONBMJmpE527EJVUzqDMFkDZPTwDRacKjj8JgIUfNxEM+ASvkdAGA/Vdo7yfExdX
LIMFA9pXJ7ZHZ7WCIGtFdssxgQlSQswIEYw5QERGeKa1gm/t7WNQ21kU0CBSqTTR
BOPrcOT0nIQiZorbCP0FAfsYokzmKxDqilmBkRuzEEl1slPWYeFBn/vmfTt8ZUSq
kgRElTweSTRV4XXRhTI0ZyFB/ezyAKoQrCt8wbP6LzI4yROvM714/b+qbeQYoTno
j9cqdwDbbyGnBFtAcvoaagmSC9NajZu3DbCqtH+SCFxJTsOoTlTBfpbhewZuw568
GxGC4rht7lj+VNcW2O8YKK0nan1hvuor8tx47uqGzCT0IKRJ6IrkSdroZOfC3MXn
qqgTruu+qn2XxERVfsZ9goJxrdWQCtWrv4l3X6s1Pn4i0C56MyXDxwQ+wY7pzOgx
4sBddVcOghP3kmK7Zp1UE/Z9jYo7oeLNUtkhFjU5JekjMyFJX7OGL2oxYYUiZKsX
fujC7bvsXE4QSwFeLW5FR9txumpu99Yy2hxOyRz25r+MvcpYFCuGABcfKMnvIzw1
kUKBOro6Or20E0XeN5wA+yUNCV8Tf1fYIZcln5CByFjzBmRl+jMFGB5MdtjJgTHi
O86dTQz95auAYYM0B0VZpgUlDGIq2LIwMTJdChiBJhxPM/tTG61jtqaGNoR6OGSY
7N5gj95I1KPQWgMCSqGIt4Fc9bfUQ0GQV+g2R+UovHHC2i80i6ChuHNFPSP/cVlN
gwUWz6gFGDl734K45PHeTsUXTteE1hH0FZLO8ET4bPGOkij4QnZRLAEFPGedrCPx
KkIV47nv+iYn8TM81WmXudcpq8fICwpC1Z8YTZbWmQTEgHGi5BMBUS2a8GmqOvzE
XIhhPu0j5FzAngH/g5zRoF53hbZ8nSN43326LPFJ9jmK78E8bd4MQGE0TPP2HPJ6
artBBEpVjof6pax8y7HE8IDkSS9iZ2I6TREZdAkY9HNR7nhLzUD6qLVXQAZ7LlGE
Wkkk12MhIis6gNpOAo+AlOR/A1eLNru/ulDI/Jha+A9JeXnw+AlxeRBMgRXaUkxa
igsc3e+OotXcmSDfmMECtimhrdcGRQajIUXr+PRdyupPfqd/PSFB1MOIQd38+/Dt
WO9nWtRJb09sJEjxuYqEEE3LJX/aoZdHndyfev5p9DrhjbqTeUi85l2g1LHtZuO/
O6XRJsrqcim81jXNemsyMCW2ibhidYNKhYCdL89Tn3P5GL9jZSnfQzmAD4Ao/hRO
uUgB1KRjOv05hi0otmbBQ8xZ1k+JQ4MOwztaiieDTq7hktI5blnx+u4AULxuB3F9
we2K+Hp8bldIyHxsVMP0zYvPgmev3hqzwAiiYwQ17zzDJEr0uv+TrLOXLFFBBPzz
/kQ5xqu/u/IVVLR8hr46gf/G5Y7dj13boa89SWOpUiiL2rd64OilAC1ljhW+xWa6
8/ftPZyjUSPvh3JHAZf53yu57bQvNexsnUuvWX+/M160tlTChyXMcy7T/9sw50wT
VjGATQVQdDSiDxw+cCgg3fev5mIB1H1DR8ywsytG1RgIwy97zZ5YRoXtknDVq9DL
k/zfw9vwiyInebLgCKI/41Jto4gqK+WbIFMC1L/tyExcy75ccIyxTqCKv2tu+m9h
i00EumE4aZIIRGJAofiKtBOHOIc8XXmRj2Sj7RwwctIsrymxTGh/5o3EQO1FyRRv
4uJcGgqQ2P0qN72HQNVUgDIBmMO/73pmnbfuYTchJjODpTAH1YyM9naIJBJMtfvl
SS2999GFsfdtwumXHVn/Y/Rna2DKsto7DZNZkn8fmU3oermZRR3tiK2R5g5p+GRG
03nw3CCkc1VpumSizOtgFhCqcCUJz57DPx2OhnlEEt1aVU4vwpLm6ahpexwqVXX6
viyv2UBjY3QBzbnPwC0YFMyhPYTBS6pNLc5eiJ7aNnffxi6AtwJiNX2QQSIK4xZS
QwvBICRxW0/EWghoE86EkfQkLAR3C1MSxjgQ29xzJ3eB0WmaXnRi1Pdxq2VfDcB5
rmKHrRUPkOMn4Ec7lowd9jSmln5LOxcW/QpD1ykUQFCoGUshllEHT1Kvn/tGgjg/
AX3NF0i/ZYckUStRL3z1q5uyI7CyPkVAuI6/IvGCThTOmZyL4wqzHcM5PnFvP2Lu
fkHs5eaysjKBn570rToKzKvWa11lCm3feAFhU7K+2AokxneI/Rxdc3e1anf90jhT
dMBAq6ub774lVr1EIdG5m/VNFsSY+bMyxoQguGmyEJ4ez3MAga/kIZFwBaXIOMSR
e9xkYa8OqitgKwfg963Iv/UJWN6hnb3EfkbntQEbsMlRR94MngS3/6Kl5nm3agj4
9+OfBdYCYHFeID3jAyzbF7l5gZe3f3/10v1H3HUgw5BC2XFdjSGAiuMgXGEZKwMU
UyY429ZSkKcJ9RNEuQlPHIFzAnvfnHqFEYp+6tIQeGPkOe/1IJ2y1Q55lHR7xbP9
ROIPm/uSgpcofX5C9vDLBWCIrfS0vWGWszrvPFn3OcZvDI0sZ7vwo/wjQBt9XLgS
e0oE2TPwjjdIIopVvheb98M+ocoJP508cKR6DbwjZHODqQYpUguiAiOmEKS0GWA8
n/HdDOLt8uW6FmpzzpZIwdc5iL1pBU5AyMWoj+bBQhC7rNLkJA+qtAsxJeajeeH4
jtLhBY4Wpc+Nf5TMVj+7WJESAgNBxeheAOBsEV81HL//8JMrK8UJRFunKYq+s9Tf
0pkEjn1YACObXTTEvd+hOjHivx+5Fm4Fzf5hJnr8R9vxlGBevPFtZhgNLW0x5LTa
5AVnKPUuY7KCOgRlyJKAWRHtyoCfF45QMZsVKOldIXCsr5kqE6PC3oZYL1qrHUDL
1PnLlHh9/l5p4kza0EJDXZYXjqZby25EaMJVfN52EnxCtQf5MhO9Ai9zcFU+4hkR
9VjqAWrEh06YQgXYKUTzx1uFV+KhOv/GmJMpJ99S8b4Iqfc0qcOse+1CpfXaZzMO
2HH4MvET2jcwQ50r47+Ts6nvMmirE7KkMztHrkWQ7Z8ia9YCInidXqLirBnfeoTS
OtHtMdT4Xv9BdOd/Cbg9IBJ60BDNvP5V6RAi1rbAlMJgje5wqMKw0EDhUbna+C81
azN3sUItULhpHLLdaoLoAEaLGvF+bTcbjPaf6AjENTo73dekKvc+oOlau72dEkJp
DeD8HjgL5FmN/YzNZtInh/PqOUxsfjyOfCv+ltDPSqrNmxCefWGTXMFfjHgxSPNH
pQDfp4nRVuPp/TPgwniYaUogADbiVnGCSzXtUspiMHWkMviU9EFJ/hi5BnxBtoMV
z/+cfRdE1NvFd6DblFFkwN9f8Ax6CVquESic4wlIf38t4lM92dX92aiykD0y0oYe
wzdPih4Me+CiGdKFmapbl4tnRhdOHv7MtHrq/qKQvflMtaxTqo1M3G8cLSmAHRWO
ugcE6m0k53QdvYll4R5MFH/gjhvIm2pI7wCd2rWGHboBth8QwM3gORmvulalxPDR
pfuec1FKqZ2GVtbW5VxRFj9KIHPTHxVgoGouPYCdAcUt4spHD3jV1yjQoeL4W5MI
2tDjgGn73ZUhWSIBbg6W0yfTurxqw4jtRzu8Lsn+AJLb1ecRZpqQ7AzFdYGbpcoH
M0hz2lJZ1Z5tWR0LqTRRvwiBXK17by4qbcNcIYeBnFylSQ9kcJbEcw4KqlygggPQ
O4VxCtVSVMe52yVWtCeN/Vf4KdXHnynq/kLyOQmqa/ZPtcDMEdnFaPN64ksfMCbg
fmuoTJOomKw94z09eQ9vFcSlHpIMeaoqxHLvpokG0ly5RVakU14F91DGWBWgF0ve
Ad7u3j5IOm0o7pxlfFmanX9U21WB2OumuR99e+NXoatk/NAkFYUnHAsGsgG6aOV2
71bcdD57j8CcdhjQta1Z5UTwVKlzzJFrCHJNlXJj2V4Jf+8nCqDuk52HGzb9RXJz
eRranNEVVH1PFgVXZspMdGRRnT+751nziSBPqcif8xSCeEPYGq3IJOtj2A3uFw5q
ZNETj7FOC+cVtjiEHiuIeUrKNUf7Sh9UrrP/3EHPKGv0j0fVZgSdrNADgFvQMP+f
F/zMszMl/M8U5ZMd7OFBod4GxrKwlmFJQiLh6pw/KOgAZ9yIMlSoDTBWbBaCdHar
jzpXny7SS7928+ZJzbydcwLhH3mKdSsaDM2RSE0qsk2Nyn7EsdJfJqFqJ8ung7uF
12Jx/W+GtQTWCJqAwq84oz5zltVFFl3lPyxR+cSBAxLy5emQfdIyRDnh8QAdl2lW
MwlCOlqJm6X4HVgwojBXZ4dIvF9od0TN4IquSvkZNdtiUCW68cRE9QCxyhnn3hZ3
ncFktFrrEOzG4+i5pGigQbEw6nOUvI/wgKm80gZu0QquzPBR78hY4++g4GJm9XTU
TntIcMcJ+B6OaN2tbJXcxeenv0jQasfQXsl+1oQvrE1BNULWJJH9BIBUqPVlRiVs
nurRPtEhHq1lg103enisSZ5e47yAsbhMs3bSJSiZUFE+CdIsR+C8P3DUTXBiuD4S
ubbfOlmkPxO6YGbOGr7cU5V+f67Y6+oA+OGzDC/vX0IfboNenWm2aNH73Dgfil2W
503hR8MuM01aMZ979oFp0jc+aYUnX5aLxeHtIJ+HDwiyLamTvujAcJvP+iDLeBcb
+ih/Hwx5jQqM7vRGc34ydRGM2sCU17y4Nvqp08C8ZsvNUZxmVq7xdjqphME1+Nn+
e6RT+Of1aMjY+zBw25pilt840vrVMygDpqONhfaZ3FKIFDOvl6m2nUrWI6kAQcO0
wuA76yKai9IKX21FiitYcnyIDyikC+MTkVo65I6F30jkTMNXX0jathqt1lAn/DGm
3XShZU1hQuCylM02FB8I+pYNADjI9EBI8so3Fcyw92tftM6F7BbyiQxz6jzZYO2N
cf+fsnnCGCiWh4xcsAbD9AXVFOlcwrL5Fq9LFSegJb5CwB9q9mJc51EINSHzhPKQ
Zfq5bkACmV5crBQHgaDEV5gjGqe4ihbYLqlw7TbkpF3icGxj8DUwx3bQZ9GPn29L
qJGeXLVkI/I170Ye/39Am4sXtlz+AKiE0SFE0oIjziiZDOuZjZIUnqdrGsZQe02m
CAsTNxiwCqrh2nztHxywuFD/ekhBOu1jy9P+S9DBAY4YnozfkbAt0KC42Mf5rwTW
X1/4K4S0o2Yx06hQf5wYYoD1X5Gzu2h3R6hBDqyLk9bE/nv3iKbfmoHuYe9G60Ks
YvZ47GKdrodjTBHresisuB0OeS7YXR200JgJ7JQU6+4p+NLX7wHcdNeLcLbi9bBV
Lg5HWCAK5PeCDvkGvIoKhCndcFFvUvDM9XdrVWhEhir7WGfGbXt3PlNkf7AqkKNg
5a+9wYLasu/Zccttah+W/V3fnrhVOG2XmuQxLRyAvwRI8ylMfhm0/sR+429mkwVs
EgnL39wo/iRaVqs1TixRRE/zh+axvF2qWJ9pbLXqRM+2Md0P4DSESWMmoPUOrpoj
Cwvrqzy4nvl9RudeTOAJHEG5m5RFVt52Ufgch0KW5Hd7khk0WJgimZNZCIWAyB2t
Lma8yE9EjA9HjG6l1CH+Zc0qWwfpozVkfHCfxXOos8qH7I44MZzrAhfxg9bq2KVh
Q/3wYY+TSUYJ1+cv1kZiumHksOEj6u636ZJ89snncSyNBkKiOTS+TjOXQ7yeopvM
83atsiGZNJDbFwj6FI5WGPteYoAMQ5JRlKbpdB9mkV+Q86PGXx0qXwyYVQggwUQD
oSMXmdvrLidUe7M94q7F0zdbve5pEgpYytXh2D+e4/j9pZgw8R/NdQ5qVTvbyruF
9Q+e8ex9TIybtQKg2Hd9KkVJvPyw/y0FZXOfl+B9UtxlztWRApRM1DjP5LI12MYp
5NmPt/6/2LQKStwnbmCGWzhOTGqdMx0MC8w7qtZPE4H+EetvlpBZt+4IrW9T8YZL
O4S+qTdZIys0XtmNnhglmfMrdkov74t49k47jQO2yfSOwwMF2I3hKm+iUwlaqXHm
0CFv5l2n94QvJ1gdBFqVQVP3EalHqhjD32tAGiqKeYotw4vM0lhpEHTjB1vtVme2
5sMWlONSPp33V6TMFIkUSDZLVQ/ue5qP4LQfMPDMB1QThAJFN82rK8njrsgw0IpN
jjxb7DIuta5ro+ytpp46G68A/DZFJr5GiN7Ty0Mb+3dH2NdqFcgz5itmRxYfT0+C
iSsr7WK9xQQu2KwvY216zGXbqFZ/mbuGWtHkfQWdt9WTKAQWzkbcx0UqB/5jzyFu
G070odap/YutrMNUwDl/bS4Xb6cSMfSM+Dv9ONLMXqZupdncceCMvWfPse6LBQkR
nplND91ocpnEHAwTc1jmATnu3AC5xv7MvmPB+roHJDKq9iPX5TMNBNfS7kmre+Qn
m3Q5hSOCTW+Co9L2EbCZ+d5pjCXbJTtabhQzNf/BW92WacMulnjEDtqXCNiRJKvu
Umw1lh6l5ODDoi/KfvJQbO79HQEKTUFn+au+AYos2jEx09xuoWSeIsvZ0pOejnpm
QesutxMBTHudlQUK2egt9BAAbP9j5ZMnp/6yB9STpe1ELJvCSclgK3yR6cd40LDy
ts66KU+pZtQywjX902KNRjV2OrfB++39KjGx1P6YYODYxeU/X0M6S9k72muQsxIR
B9/IEoZmmnpK/MGXKHzxnCyt9KecyEUF/IOIUlmMGfDWSrwi1R19+s3Wf9H3wxdD
XxxVe1VrD0wfUhCxEUSV3k4EqrNWIvkkrPogLBM3B6mO0gACoa8ilm9aFySzHV6b
C/jPyUfe3vs+LGgzN1IPHKeGeJfyxNV4IHukjRSh6RzOqCW7rT9Wir+HFXGHhsYt
nWXaXKoMUMYNsH2Tq2+k5wJKfdjzWP0gAijwS6vgxV5MlOEtFLOnvgaAiDPDu5o0
TzA67KI5R+R4jeq03ZnHDIleaNvIB08yI3yGebqzxafwsR4d2HvGj7MGSyRHzp8v
Q8qyhbeg93ZJcFzu71SAlfEwtc8/YMBc0bH/Ot3puUzs/B3vKZcG1Y7ZKkQVYWK9
yEn68809bhjChhodn2eIEz20CUUPrXorflPAgLhCWIifNMM2dRjNsiuMYkrIj/Yw
fD6m29NZUxgvA66FcppVcgYOBUhSKCK6nnU4m5WKOuh1cWwiBdXbMwvOv16WoGFR
qWgWcv6w/D/gHGWW5qryyFp0gvEvtt1K8w6yIU/wfNHbRKfuCcPHiuhiIwC8G0vQ
nhzOAuMc18VEInEZt55+laNklSO4pY9CNkHSP2tp9kJ6e6Gv01HOpNsBTjXx0lwM
F4Bn3XJDTx+PEDIbqZJ7FDACLkQA+AoLl+jKxd0K6lv7qkjzYMVKwKr14weIxpPc
HkbX0RU5nSuztCsgdckyvq61FjxOrxJr2kQUZ2ptaCpnFMDtCDPF9kRFfQlT+p5F
UEXfLMe2cxu0tGRvS94i89szyUiwD3UWe++J56RUOp//AXm34qPgYg4i/4NEGhfa
uoJg/4qvR+9BH+Ay7/nzxR1zHREj7dp7dzzdmkeFn8fPRxQazGK5SLKtKO93AIVu
A2BZdcKE7uliubBAo7jw8iQkyenU8V5YoMcU3RcJWAB0FKVwaAsENc25FPrS1x51
E3P9+6G8C1GwZl8b5rBTS9jW2kURtMeSrMWoBAZTvFGC+jtWPGfCK3Gtowmly+Ko
mdzbf8Y730rzhAVoFcYIhNry65gd1rkL0wmWDlEY1vmWO9zpG1esbEhIOTJsepTJ
NBJ61E7eneuCiZAtVssdS0xaUiHZvfs+mK1bzMeOZEt+6tlh3Vi/4cROMDMnz4nZ
4Y8Em0lTq5txZMb3ks0tlelPvj61xAjV6WjNlBGSPZ0Zvn5i+InCfb1xQV6wpksD
frN+aZ8sB3Vxzdcriwa0a/Xeao6FVpeU/+par0f7uoSc8VGKWLPQmxEWWmVfaXIp
o9N6S5O54bNCzEXBY8yLud52wiLxafZNGDwyTgkTPO2LNSb5c30rGb7RTb9+xIDb
l4XdCYiKnPe0Ex9J1T4G4Zpq50dNsnMW4YVAXZvIURoG5j01pXvTh0UQI0sOM8Bf
FtyJCp579ASMwi/JpFLsjmGE23ia736nR6Bk2RKW3fxih/RMP77d5LZT6hMjtONK
Wygy+wAFGyqy/7fbNLqvye7oAAh+lrtJyRqOC2c659ibikSNFgM74A6+wdTNDqzp
wulakMvbXNv1xqGM2w8dWR3ioMMTdOUxm08xWCtf/htGPPtscdSbfflK4ogk2xBB
LQkePAd7wRz+c0mJuIxHj6WTLPDq5oRK61XBeZBwLwkHvD/ZviXK46h4wavsX7QF
3qmUl2hgEGZ90Wh521jiVzZ5c8EJTPKpg3KXjz4sl4NtAMR/dTVf+eDX89mYLSN6
BP55WaQIiLx2OkcRdJhbESArJBlvVdlCjCzh1Z31YHrCuytxRaQs2P1cQqt2j1xt
Jlq3pgAX6bPNBOThaCpl0XW6yalOauXIJRsvHEXFK94aJ8egtTWkLUvpRmzLpR7v
bfoQ5WEQTZpqDT7OHgWfU+PJBGML+KwOrsafRPUMGoIaLGNKu8H4oPAkpdmV+mzn
y2zGWoGphutJBGEW/1Mf1RH80U6s56Tf2L8X81q/qSjqaUPC2ipNaLgIEyE706QU
OfK35kmXGI/e6jex0jbX5j7ZeOkmazcKkBukpTNmlqYiOEJ2E29prT8eLqXNvDcg
OehUjBZPYqhSVgRPZf3RL/YAyTl97N8GVfw3Ee3u/4z78FNyYozPNyB1JCRQjIao
AoiutBR5ioYbkJDelMqdBO5xH49I42yvfN4GM7XUV6tYtbov7on/AOpHDc+40x5w
PS3261U0SXM0m8bvn1P9NnNe+4Drg0Ij/xCWlun2ceuRoXXyudxT8CLkDepvMXor
jBGzSGWZR2LSehb6J7oTTFTNHl7Ko4DNrZ7t/KgbO7aJ6QSWMuTQ8HYeycA1pLfH
WzWg/FBOf57z4cRFm6hsut5CO8kFgvbdCtEFek+qQ/wcLrhS1chTP+4bnaw8UAOd
W2C3m2+zlMImQqLmSjy3qBeDRS21mOMq8uiZyT5EzoVSLcGhW6HaWkd7kj+VoEOL
f9zxIAepQKXkr3L190IUEQscQmX5a7wa8IcNsnM9RdFnDRVZvNYiU81ZDNzohhI1
1w27XgpS/yYhMyGDNO3Ab3pmcwUy8D8qu/VckB8TfiOAo4J1XP9fZ3BRapCmlK0N
EFsMUAm1IXDv3EuLw+Dq9Q5JxPbkVkKZs+1IHMGtNC/epygRORavx+LDPG3IL5xA
rGeWpBdKJJuB6c7Vn9X33tc7k7CmgOPTGZVc7igiqxQcTkWwbAbLL7/RvHYldpKN
0bKEoCxh19PwWAZ10TaoY5A4PObn5c/1PIJFDFa+8mRMe5K0i6nkD9suaW2M+A6i
Y3u6QNmPm7OkWlDoh60MX/WI3+7XeKiyV9OsPf1hOf27AQ3mZm6U3d2I2EJzuo1B
qveVrgjvavRBETb+lfIoTq327i7m4+PA55FRKnlTRbbyFslLCfow2k7Iy/ftSIxZ
Aql5aVjrY/PBNKaFzQzTLHCSJRYBnwGk3tJMZAn8rJ4vZ1S7HEbF6p7/dq7dyM68
Zr0InQd3/PEUM5seqJ/dkM68++euO7Mkprht/ZQlMQ3pnGo5ykqNLeU1hiGjtr2c
M5B7QgweswusPC1tbqc8eJRDT91RvObcNLTnjSCF2SP75ZXmlIMlUj4SPO1mmh1r
aCw59Yv01ozZrtRRy3dGDCASyRy8qtNgpBSzHwsQK0IiB7GNzupJNHIcyvCgyN4v
XSqvfPk93+JGLHTx2ukh19RgAOVFpPMkawK56HllwxzLdy/Qsx2ODYe/QeFDTHX0
1iIAp7YFXOObmGOafu9Grp5XLWV5llEGzVKxCMIyypnvpy6amUwPnnycKZE4mVsx
rflF0t4TRxYQLq48qf7VhD61jOk+d6DtM+su3cxWKsISlVKQN+lJo4rraEw8Hx5Z
bzkGg+GFsHwphpyqqiEc+Xi0l2wiVnp3LpeREaZfHfTKAFLG2YZmlYf0Ejo5ddgF
tUPoeY49OHwODfaWdPWcW+xEZlJj2QJcV/wSFXFzXk+e2Gjuc2xPW48UnCzGH3bX
+e/ZaCkrMVmhs/NcKPruL/jwzxVe/2KOtr7Zey41tn+BkovTtPf+dlcNVygZ4m8u
vqLKAymmag3AjD4EP8somZO5v071fRiBCB6GIl0NOuTCVoDm/5y6pSME55p3Ta9X
izTRL6MgjYlzFp4PlAhyiijTWX2xQPbuQq62/LNj7QhymPVXAUYyc7FELwIVBom7
mkQMlgYDZhHfEBjpN/75KaFmoGuP1fPTeOSTbzCinMMjD+49wFKn3tIVp/j7Vacb
0PtosbKyH5946HsiMVDjvZ7G2hD+f9wc2QfMj2lQIfe8PoY5z9IzKERwahBN1O6k
PGmSVn+U3cNE5vBlhzBUfJ7XoCNYps/j+MQVfupCL/hyBSZcHPkMlyN97UoidrzR
jiOHFNKBXo/2nB8vlBVI/Htx4V7FjWIyQ+bmLKbya0A1l24hwyIlgB++A9uO+ska
V+VVzKwtXnKYZYT/lHkSxTDoZuM0YmKIWDvlBhFq1wO3XdWI+DUVgHm/dETvHsiK
EOvLjIEGDiAOCsRRhbQnBYsDe/1deBzgo7Z4pFEL08o45QLsFLrhmkai+D80Nl9N
xMPjIJmxAFuxXhJKLMmvTGhwxfM0xc5TwSsR68ZfQfKDWlgwgqC0rJFcNs5Kqu5z
7rXrZ1ZyCPa61A1QDey/yuI9xU81j1D6Brdy5dHNJuf+iuSdvsYeqUdUWRpaVJeR
up5fxK2baB6UBD42Q1N+vcy5RJM6fVr7e0EJkNV85gCsHcJTVVHo+AC4dWYXLtOj
`pragma protect end_protected
