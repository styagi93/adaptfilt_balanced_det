��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[<.[tӒÓgx���)1��i+�K�SY���'o�yM6�`kNX�
���{A����R��%�=4��o�2�ИD��ȓ�}��t�z�-7yD���)C��<�f��qF����e��I���8�	v��(��z��{��WN�'Z��w��&΁�R�~�%��Hp����U�/R+f>"rE�;a�=�_��k��L���GEnfF�B�y�1/3��ro���1"��� Q6�B�e��*|&�<�%�7o��(f�m��_��Fr��;*��y���ڪ�f���$���%�q�K��4>�>j���Y�#馞�hb˗BX����WE��y���32Nq45﹈��Ir��Μ���c^M.�����V��?bd�Ys����=������P&�Ppj�c���IO����?{Da�$�-Z�� �m�h[�n[��!�ۆ���c�2�<�-I>��3V\�,$w��<��@�#m�n2NF̾N���d7 >7HV���a�co��j�*�*�-Y����	��-�}�]N���Z�g�H;H2A�es���n,|�$�R"�ǉ�
��J�Q��p'�α�I͈�w��6��܌"W��I��U@w�	BH��;�~����8��ȹA51C$�F�4$
�,��<)o�~��nf�`��%:�Q����}��ip���UR;���F���0���J�Y��o�J����F!@�L��B+r���~�DC�o���f�f������{/u�G�DIE�ۮ{Y@�CSZ�JoF*?M��:������6\_6����¤G�[L���a�Ux��L�#�f�@'��PZ�V��I���1���M��*�ɯ�-_g�.���E�O0���~��I��|cR��/��|�qQ +;a����*+n���� �DL�Y͎҅�T,3���c��we`jRh�B�^< ;��І��[WJ~X�%��d6�8Q������1�Q�IzU�U��͌��;F�p�oS��o�8d�yN�����Ǽ������Cx�2,��t�T�ֶ��ǳVH�w.��ة��_n��&�0Y�w�>6��៦DJ���_I8c���]����1����L�<9_XtL ��̘5� ��8����^�2�֡�`�j���z����b#Ζ�4)	�7�����ԫ�e���^�^;L�X�g�%(En�Q�2&1�?�W!,��B�ʛ�5��h���f�\c܂V˫��]��{��N��+������#YKi�����)�Q6�u~�Aڸ�&@.�� _�'�b.Ϗo�eo�4)�����l�^k@3�'%�tͱ*6����R�����[��[�~�J�g�*%̠�G=���{AG@��9�m����W����m�|ۺ�ѡ*=�}�UW���J;q��:���]�<R��p������J~FW�H�7EF���&�pmg��_49Xd\{�*�I`Ғ�z�N�Pa�u��j��1�j���C�B�>�t�ȇ[�а�	�7����ojp)"ȰutC �n^�+&	W�����L�C<�����a��1��:�,>�!�m�(�ly8���V�Z�3cAy�!}G({���ЖX`"��V��M���αٞ�b꽙2S���\����9�9
����\j0DQ�-����b3��1\�)�r�BP�w>&��]*��J���[���J[j���,�dor��C`9�D�|�𯂰 4]j	�����xQ�H�qĲސ��II���U�y�	Ҁ�Ԡ��n�ٸc��߄�n�*Տ�7�QW�BF�@��Ԗg�m&Q�|(�N���>�{)��y/�����m��;br��GY��rZ��w��^K��d��ia�2�D��vD�^�;�2U��w�	�"�GRZ���Ӆl�pNdi���{�x�vR�l�C4"�X}��lN�&l�z��<�g�+�֓�J�ɥAM�M��:��4�����gO +ț�o�T����sҮKF�^��
�Ĥ�]P��{�o�n��-��"����_z;�M�_���P�y0\Q���ö~�ש���3��|�G\�sЅ{]B5��&�g_���gLG��
/�fua��ʲ-u�݆�C���q�z�� ���	��n��h�N_�����d��V0s���综V;��z��+��!�լ>L8wؗ<)Q?����8�yMP�qʆ����N��X��-z?�ьc��З��&ʝ�Ba�U��5ė�&�'^�
 �
�z8cC)�� QdԸ�S<JT�޹v\C��Uc�M���Xgƨ(��@d������B[��^72�i�
f�/�^?~�.�����_e�о;@��s���B�S�`���L�)�b��N�;�5��|G�q��,O����� !�\���.W ��(�ƴ`�(5Ĺu��*�Ӧ���6�3woU�o��3 i���x����JO'|z�S/��B�;�*����Q��?�(-B�A4�X2(���C۽6hU.�T葪`��������n�k4?N����0���I��wa�w�{y尘��M]���J����{o��ZH�=A�Gy�@^�B�6��K/�j7O���5>A�X>�,Yw�c0Q$��*g���t8`����-�:�~L�v��(�T�^H�J�3�b���� ֑��w���=h�qB�ĭ��a�:=�@�}�0�'f�6�G�sLe �bj�#�8A�;<�����O�?�����Drya�d�t\�_͊wn�̤�(�����HB�z�@Κj���`��2��#br�� bK2�WL��Їx+��M��A��LW�,P
�a,�X#��$���6@�������b*��-ut���k�y�
r�M�޼:��	{tT�����[ �7�m�L���_��kn��P�=	�4c0>/b�.Q���o5�֔5���ڂnY=��
�g7��-��Ҩ��� �쫹�]�=B�=�Y�pNm�T��Q�?j��H�/̙)l3E��$�NY�f�.�1���ii��>Z)���v/�*�խ:Q�&hS�K�Hb�pٰ�U<6~�j}?�8�L��� NY�\k�}�&k�m=�r��Ȳ�x�|��t�Ϝ�jp�)���xS�7�-�$i��0��h�5_1�쨹�)�7��cB��"P�u�%��X}ҹN�+<ܠ��5�\N���8�@��s�/g�s.R�nVE��P>��F?��W_7��
%��6�_Z���V�$W��	Ϙz=|�~�T?-w5��X��w����H�#	8#ε�X{�Er�`�%x����^��s����0F�gC�_��ȫ�Nȵx�jn��8r�������6�5��}c�(,:%�T��%b�D�Q����ǂ����d���W�{.�Å��L#'��&�_���K�b<s9����.��e���)��fg)%b�&��a��V cUz(Y{�5m:����.���=�ïҪ���{��m/$x�)�΀��w��	�A�6I�V�S��UpR�2W�zS1��z1G h�
$��C�;t1JZ],T<�g����y ��rS�90�9��xC�R ?�꾤�o����N�d�YK����~�p�R)�AV�:\\1]�Da	{��DyLd��2It��\>eӌF��G��k��U��7���{j��u�XF�Ɋ�8�tP�mm�4�~V�4ɡ���)=���b&E�a�_'��.Gu��R����W&?%��D-���+�
��rG��R��U�!_񑻷���sY�q��{pb��]zˌeꝌ���E�iR��
��>��׃��[��7�� 7uH�[�n��������ۤ(巿��k!*�Np�b��/Q�p$���}x���V>���`�-g�#�#@a�EU"�Ѵ�ƻ��k#�R��0�T�?��S��5!R0���>6���v"�P����Q��01d��1�!���r���1�ʝ�.ȳ��G���P�Vl4��sI�)��	E)�n��c}(%m}��W\�.��iP�3��+�{�:}���xf�6C)�k�(7�}�%3�e�S��_��w���*46�rЮ��Fz��Oy��<�*��ϟ�@���ISu|�x� �$��b5GgѶes϶$H���>����޷#?��)�.*�^5����CE�0[�1��m2,尲3S�4�r���w���o�2JsX$�3>c�N�{<(��%с�cWnAŹ>�g�e93#�ȈR�3P�ƙ�� 08X��m��|�/1Wk�Q��A�u/���҉e�V.2UA�ٚ����ZG�	W��3�.I�L��8�R`�r�^����!�9�] -�:������L+Y6�`B�P�B6���<���?L4�@[��U������L� ��@��;�{OU�}���;M������Ȑu`e�'S�[Xj`+��o��y�/#��e����wl�����|u�)	:��/<o�v�V���WepWVx��⻍��L/b��n��lw&�O:t��d�9�r'J �i�a���ܝ�xZ��k��V1:䅴xf�uͫ�w�� �/I蓴���?�li˂���3!�RX�Nn��f��^wb܇L�=G8њv���}#3{N�A�9H4��ԯl�m�C�5��5�&<yl�%�p2�x�ܑ�wl2"�N�����CV1�#�}	�����@e�� �
����"�E�̊r��n}��}�U4��Q$SX#�r�~Ʒ��n����*Ѐ�!��c}��8���7ƇZ�Ό׮�W
U��W�2Dia�!��2��	�5LD$fl����ae���ȭT�@�%G�h�'v��w�����c'�C��uJ�(�x+�j����4�6������v���K:�O����g�	[����׀q��>(�aMb�d��6b�Rk�e����r9�/��Qw^&y���:x&Z5���#�~{%6�O��S���t�B�&M+h���p��4�Џȹ{wK|��5���i(���s)>���Ƙ�i`�3��
���S%�Dr�*[�R͟4tJ�:V�2�Z����zm���Fh��Z���&:E)';�g����7.�����:E�B�Ds�22.��}�^߯�5}㿷��R���!�|�n�����Uu��ύ�_�盖q�=��e#�rҁ]�]�Go�7��;ƫ�i>�P� ����I}�� 3%�)�������JDizǲ� ��s�>�e?�e8q�o��Nk7�2��f�s�p�"1ѯ95���a���Nb�}a��-�P��Ks"���_�C
	�[�t�v����T�^��V���Y�UB+�G�h�5D+��x$�`��?�Sz��:A�U �ȑhz��%Wh�4H#SQ�����1}��b�&�j�>�ti<�Cw� ҂��ہ2>"ER��	�^9��M�zEA�:�����VY8���k���R@���|?��Й��wE�#�R��NT�xk�2�0��`s��Hɔ^��	0���|�zO�M5����^�_���2y���T1���� ���:�٨�Om��6����v�8rK>�7�v�� �"-A6��ˌ�ΠR���xڬǘ9��7�������
�SJB��aR�3��S��t ��X-�?$i�J[MCp����;m	�>�����b�ʬ\P���\��I\uzm�z�*
��q�T��>�\H1]�K��s�#��L,+�F[	m��?7��d�T�>0#(]{剋��;W<��h�4����/5�����}�`����k8�[�G���&���b�i�J���V����{���yY]���}�M���O�^H�.ث�Yr 2'��L��J�0��Ƹ�`iFY��3;m�,��#�^g+r�RSln$�u*�HQ�F��m&�{M�.��p��c�o��A������7��]X�)_���p�r��P����#�Z���F�,�`
�rE�l�ǣ���v�d0W����}���'s��?�&�b��>ژ`��@�V�)f�M�"Z�&�tvb� L��_��=�&aХE3z�"���H,�D�D�n��K<���fq��hu4 �9������u�$	6o����)��\Y �k��s;�6�+KJEd�R�%�w2�g���d���˗�Jd�J��G],~ !�S�����,�Q%'�X��߷��6����u�VV  ��G@coL��ߏ6[��ʦ]���3*v����<ߙ�d��Hox#�l��UT]���D[䰼.��Ž��b�T&���D��Rh+�SJ1�}/��QQ
Pk�_���������u�Ϫ���z:U��vO����!o����H����1@ Q}JiRat[	X�Q�l��fK��j�������~�$aܶ�@?�"zA.%�c���W�����~��{��D��
�D|N��ʨ��mkx����؀�J�&	Q�Y��dZߕ�L<n�
�v1o��^������T~��݈17���Ec@�B�Dmd �����+-U넁������� N���:���lO{"J+)�Qy�c�硍����Al��!Ȼ�EC�ov�1���������� _��\��T�ć�a��]ܔ�\�?I��v�٣�TY���W�{v>؟HY}f����;J"&���4)��`m�r�S�7�ՇP�"�3/����"󡐆M���N�O������Cp�$B���6 ��0=M�3	U�����^C��OK�:"��i��K��/����]�F P��D^�5��W�P鴮?J���y �yB<$ux�����n|��گt��J����ƔX��Ruw��
�Q����*����2����;�����1����@vm��A���3����3�+nM�}��z�D��s����7��x���@k����X���_w R�#��W���v:��!H�j�6�*&~�U]+^�2: ����P%�Ռ)a-šSXC�W!	U��(hޚ�z��/�/���=ʹ�:�X�ˎc�Ϣ�_?��<Ia���^��'�h���ZC�A�[x�� "���Ԝ +�����W�&��[ԋ�x�+գ��*��A5$��s���7����!�yom��ݍ�7ٌ�
�r��)e�6�=\�R�n�k����3����P�I��/�.ʢ���Oer�5��7�'�i3��V#=Cm�;[��C(��otq
æ}���|,��2���=��N��[���&^ԟ�8��,+{B�;�ͧG�e��]�"�Լ%�逥N�dUPr�C��씥W6;�#�}�4����*x� Puad��E.;�{}2E�n�f7� �[`u�A]ͩ�~��:�4����3�1���9yL�{�/j�����߂5������� ��߬(�ԼҒ��+�~#Z��$+�ŕ��qx^�46��=!MD�is�Ȱ6�3� j-�����~A�����:
��e)�EVcM��6�Y�m����v%�I�U`����W�s����I�b��Ѯ�������uS�z3+g�t2�Ǫ͐�v��'�6;��c���W��݉6��(o8�'a�@��,�����ܥ��?b�w�!�1�����8�/q�=�D�����N�旄��G}hdȩ �ʷ��Z%�,����	���xA)D����n����'p�D/�����ptg�C�'��b��8��g[�=��]7��/_'���ʁ�/e=j���?qZ�c��nY2hy(�{)��T��D.��$o��6d)w��HP�>�][��$�
-�l�Q��������D�5���;_����jQ���cܷrK���~Y<q/��y���>�ޭ��·�p#���73`����k���V�
w�N��\>ݢ� ؗ8��-f�-�瘎�Չ������E�Ygf�%�����Y<|�o[W��Ն��|�H�JJ.�(#�+Z�����