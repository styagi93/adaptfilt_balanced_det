// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
fAC5clpjwFj3wNSEVHmyEM2fEf9ewg5gQJGqEbOMePkuN4LNTXbKFcpgkcY9WJ5uaGkRNJlB8tX5
yE/ozsDZURbPkz/4Ukt6wI8Kp3c0XDkl6gvDA2YDdPU9i0/UwyaK3YePK/eFnxRKgkINH6jcXv5a
Al4umFa5CCDPDP9pQBRGZItT3o3PJ6Inyu3dwdzHfIqgsFGKcLke0LqoiyWasizIS8x4ewiP4I+D
jCMXglt0Qjp7eGAdljbUH+T7IIkObdja8UHvWn7TuN+Nhhmi3gIa4anySoEidCUuD4FGZtb0EfHV
nRljPx/HWPZIPmJv3Dm04CbgydXqBLKcuAN4qw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14016)
s6JnlsQn70EY6ey7/auarfqZKir4LP8k01iITSw+HvuW2K5RZbevDAiP4ZeJ3gM9TS789QZ+lUna
OJUt9MgKsBjmYZQY0j3zMlqNXWELJqIg7B9Uj/d+mPKOKm4sBbuJiQJn0Ot2vopfHtb59LMxT1J1
tEl0hMezSp4BWczwaf43GeCj49xQpFBIoMk51LDLQ7tdz03/c8TbQvlmmVjIx4WsDIiRkfTMX3Ek
PkKnMxNuy6SzO1Xbf7Yr5HJ3jbrp4ImyomC30Gq/9bVLNKyilZzD4hL4QrsaHhSD1cVniGl9tnUs
T3uWS9HJfKq4Hp4+TKbL85VuE/pQ4ZnbwIt8evqS5ERrhzLBngFljSaVxoyXImTKL3OpDyfeQk8h
iS9U6u87PYhdQAQFy8elo7NygAqEAOs9sq5xQTbAsnoaoHb3xcOAAEPCayQVJUtCMmGdn4NXuRvK
L+hoU/N5pEV7Coi7T84e/egt5CgxGZZ63v2qp5N5IXbQSluuW+9DIasdbnpIt6WAb1XoxsIBYnCA
P69jhPAJvsvPt81uvPCy4S8FxSHAw3/eFsAlFP0IrdW2JfooXjLK5j9hb0NyausTKGV/4MDdN58v
tWSkuK6eA3OkHsCDKYHaP5y1irmOZR3z3sVitdYbiNapEYTt7oHm3fOm1PQReB96oNQ3xckzapTb
Hhj31yc859YcAyU0XARo598mSaAQVLg42izshfJO9PFDabl0Tyxzl4nGyK296/FRWtZnFuRrPkrU
U3myzyiHiwFPa6rwYgLBI1jBPgsK8yiN5yWdIs61wNknCfIx7c7rC+7lEy9IISGEgeHbQYHjvfrY
mBC4fqRP5w/FLqf0SD3uIeIpYB6jHQyGOCzhPDedEdQg+6dhT+We+wKErjIwZKjXhrvSp8Bjy+OJ
KlNQy0CHqtPjymDFHpo2XxkeMJ+AI/Nw5u+kchQZvSY6qTcsLgdNTAjr4Q7O+35FOHtWSQcHA7+5
Gh7Oiuevlz8Z2fbpYGg/iIgcBgBJXzeWOmwzI3LGp51nmn4QcGG86DL5pNpQOZH7JKyrjg6Rr0+x
6h76gsGe0uSl61KPMhWvaXbJ7Au9lHh91yml6mzCMNFIcgZNkXNp7VUHCgSIC6FRZzGVWwjdr9IT
lRIzQlCHDMF1ahA1iImy0JuKGiBOfUb2DXlFRAMGQ9vKu4vla+BF52uGl0WYe7aryTI6ZqJYeaqz
RxXFYshbJT1CeLu08bpDNbnRnxSakfuqxD5aLsO6iNvDKYCiFvrfxqRhZCWar08ayoD6V97NwxVx
o7t/wMOIU0F9CWDxWQpCHuDMpr1IEolPWzqFPius3p7r5t4qjxJjTkgu9Baj14ec3Cg4rcuzQPel
OcbVe6YedVkSRvVDDvOmSbi7XCd1WMGl1fm24VtRKYYOpqO8bGC8cvTKiutsEMMZthfFEy+uyxmE
S1mpMF3cWOHcNU43T0lbBM/GNmK/jqFKu0VGLFZmrGOs8DTUT8INI8yRXcK/LQA52c3uFMZ2DST/
mGWscFUAfllNJh5anht4sSbRBh31rxm85TvOeafDgwGN/J+eceDQa/GMc3M9m4wQYwRFduAAxB+Y
yQm7xFmrjEQmGFd+C0PybyrViaskKehDFf95INLMpheSdVB6q2i51KeWLx3kbYGsTghMs1iX9TJT
0rVtPKL9QvzVqUpRWZX2jCYX7X7vBuuD1Tb2rlLq/tx+eLwqPNQ996ZbslicAcWRsXOzK0W3SMHQ
lg5aVzqkoraypaHy0yMRxJKkDCVp06ZGWSODrkiBY3FfnxbLyZsvDewZ8+Y/2caUp3Q2Ufq1B0Vo
deb17BAsytjNmR4SXqL2S8whRQpjC2djw2tQRwmvbxL/rHNv4rlFJrQsb/gR+i8bvoJV63vKZ+1/
D8mJynPlNPBlE5fMSg2+4pR3+yfcMrVcAalx/P+5EUFKW5tXwmhBudDx5oazYTtjGC+Q0OP8v0xf
AJV3espzbkCZTP3OZ5nWlV7pq6ySZPJ7Byi22UnzkM/yYz9boZeh4nfmNxpMJlcHtRfZciECe8yC
0qiztwQdiZeqzWpgQOIC5gM/QIbhgo9wvgZNNSYOKn9bT91pKgmIQmtBLVgFHIS0HS7Nz+Gyrgfs
TgW/2XkT/bf8aMSglRN+2UrXdc6DdteRARHAjOCUTqmDZKn1B/hQ5I03CNpRrUmggQo9Tpfv4DPX
IVlqpyRJ8g0uqnfZBSoCvoveE/qHqG90YNwGA9jHzeyKw5LRtAsq63VshWegOpJJzE9xhmKQ8wRR
4cqMT+2tBFDhh4BH26JeTKgRBG7ou+EfE7DZY4DzsMWk2uTfhUCicSU9jF2iNNTsUPY0GoX8wh52
UEGiiLow+HxD2jehLFDAN2/6FPHa8cPpCHG47l/1CsoP2RVHzxtRhhk1tR2MI/hjR7I9UbxIYYcN
E1LNF92kIhoZcBsZo8FFQtTMB0vfUbGnt/0J9+YG4nVCOkY/4M8yldPgfeQsOcqZVNJMjXd2nc1m
6JqEaCrp2MCykz9iNCeVZQDXIRpzMcDYa3tYwPj2y1AIu6mnGxpR0jM8zAwfXPKiAVVcX6QZz4A5
3Tqf3x/QEC5y/o5lNN85iINtoVpJvvc3Tr7FlLlLpW9rigLfKZBfHjaBZO4R9WZneFguw358b4h3
j4+z5W4tQDScf6FUw8pYTu7f79RZuMFez355mi7BncMIRDVZRe6czK5LiD0np3MEKO1Gm5XxU2H4
HItqYh6ZTuazH2yeiEObUSxl3ctKSV94uXBXVtXb9luppdcTj+d2oamBt0q2OriMxldfiMOqSNw3
aHMLcHm1tA5w5UPD/F1U6uB97Kw1CQaeDDlJquAUIGyIrUILALlPm/jdbSLZCdifnmPPzKenHyRn
o2/l4Th9i1RNjURxI6zpYjWLl0pcmvn7MR5EB8s09pf9VA9NrPa3XhCQCvz/EH5W8ouWBwjFYHdZ
1fiTfRdEvU3iiqt3BC3muTzYeyZp8MJmjEsOKKeD5mol8HcRWWfS+KJcGAgKH7gGB71gW1UBMxIj
/RM2kuree1w+iPpQOO6EzUSBaD97eywJuZRyfygf9NbEYsDc3EmZhtvRon7mE+zfPBri6NtN79mx
KT9RdC6qfa+lfn0TJtUFo0hxsox4gMMAb6v3Pu7fYsXLGEr3yHMV0gG9OLUMmJZu3XRG9bQ9KSxo
g15Scum+kDrxXh5nr/Ga06wUR+ivpjiGvyGcrxxWfC/Kj8gYG+aW0wftjSM9dD6NMWmhSW52v4rf
TDhxkfX2VDc5ExPpUp0VXB0nNva+IRzovrs7jTeHCe2cA/UH5mWwxd9qliHMh+GAaD80YNfEk3We
G02aUZZ4LENwZppJzTywrIU2tiZIX2NCkH04gNCNdKGQNH0gDGDxf0vknP3Bk+Iw328FoCDBHJew
9lABN5vZwNutStnimSIIKWIZXZU4miZ5uFkpmiX+mQXbclmcfmU1tY+aRlT6SSdQT++Cr2RGY44L
1b7nSd5PMmpcuq+MI0kfNw0BgBTd0/peDvEQIskxlGM19etJKzr+zaIiqogkHtPhafduyfXSLz6h
R0WUB/74jeRtu+jhkjKhKc8zMQ+LvcPgY5Ra5Bcw2vEKSHpxs349DbLcXuYly99atLTG6G0QpLJT
7p7P8tl3/O9/sQCEzcUR9NarPWeL+nJoN4zXER9ac8jtyi/iXL4P3LWiF/b7O9DF5cV44P1c9/ZY
VunVmVEtm3C44qivnfaxgIkc8vXq7jpCXDm6Brrj1bTLHvUWhDqGKNR3Fdw///X9VgVKdkGVvVc6
K2V+6Z9bSKKa3Oca4eFpqpJ5Goc5HasAvo037u+7ANu6OUWChigxyC+0henXhCFP7uC7oFf0MEXQ
UfZ9r84e2s+VSybrRZ9JBKZtU09GGTgMHJpx3t9HMB1vjb1nJ8steKNpFb/SiIHtT2Avu3PsGXRb
a/1HzLqJoWog+6YDJAQ+Q68APzkfDPN0vvzu3GATQkP4haU+c3a+M+yb9DMlcxfTyVbLk0QBsKtl
HOPDVLq5vpWljwz39fodZCccwLDMQCYxJHXmROJmkiitx2xgt8f57lzLQLgMX2SUD88/UYbPQBKw
0xjPjZaSu6vi/+0ykDBlPA/HkSG6DGJsn1Y7m1D7aU5uxhR/jPlq2qwqm1+5tFkK5UjkNx0VBzMJ
M8XpuMAbxFqB0IL5hsjmUf7+YrVQF9xFizDuevMEU/9326ab7lh3AzxYwTY4pghdhqG6gcs/O/jE
lnKRfgeG5JrgShXCUljtdOBDPzI+UsICMHTnMxGScb1XPL7GOGgw9fEPO+6hn06eHS3KIAGm1GWZ
kcI6kc1+KfURCHEMO7PI7p2Vz8pygqdoNSPe6+J2VjFpsEgk7rM1LywEWlSXRnb1p5f0MPGlx27O
AuX8fdv+VOnIpXyYJ5URVqsyXk0Qb70wpfvR1ozU5/F8mA3Ee5SwlJmQmeoUuke+kFeGTZFRXwWN
Uwkpr3zE9foYRvra4DRSpxVgfaGYUdzFYFfzSsRp2ufiZAjGCX3fUg6dzPzp7kJ0kHKQnSR5HiMY
XwjiuUtewvWB0KZhQlWNYGexosoIhCm3FUnTkToHq140JFgrIoJziD5i1zZ6lCB4rML6iOHfjKu4
ZrW5kq4JceaUn5KI4lAGmVEyXKOEtGzNmd4FpsbmWS6tat/9VhnMwwdRvcNCsFkT/3i4S5IbfgP7
OFpQdywLjcuiX6LrChCO28rvtnTOPh5NpBxJcL35bTfE6noyXdV7/EthubEDmXP3+5AgRcekcQoS
Q58Ayj3g48MAVdJznGoVIttHRrzXzQ0AaijQCjQDiwXJg+yCnGQp2JaNUdSHG3KiHMNlkV3fyCEi
qZkrHD7vf0XdzyFeGHgtgsVVYVQhDColxfCTi/ljhrATYgbV+NUivPbPZYUVAPKBaq1Tih7KuxUe
j3+C22PwvTpLq+vl+9hYnfsqPXe/6NBw9jmDYrPfaUEnMZgWEVQW64WlLSKQ5YmODGWaCGudW4Xa
ylvBgr6WPjD3iR9GDyGP+OrkzgPVtdbOUL8dZvolKvUzBpFZWTNQDyLaTm282NiNOTQPaNsXcz/+
wO2V0JEsV480DgArz/T2zVA4YIcWASBTbG6Ff9KZ3hI0SQrACd7/QAR5CsZezXbv71AQZRETteEQ
EFSz07hSj+nQntEgzxiL4A1JxglIgeq3NYMc9IX86MhVG4nCvI2uXJjp7MdXlbkrEkzFodW+6u1W
4OdTDc8x/aiAjM5LgzpJVxXjD/8a2In2+YKGPqUGFA0mU/I6hEil7GtL4DKONCs9HD3Dho1pXkK0
eibUUq5tTK3jHDOzhBVbRvEJX4WkcWaCCZMHox7G4hSSpgSQ3GEcWTa/oA6EevdgmFfl6Q5i4uFk
inyS0WzwoouIV+McTgi3r8cSoTADxAcdPrLApEW6BFg7zv9L1pEWH9k83N5s46EWOH4sgN4sCspF
/WJMiVd2EsbfX2szr4zWv7OQ3tQ5TCLQ0YdhdVIYjvQP9aOHwiVkIjTrEWbzr0x1/TY9zSW3aHd2
kKjmonu8n4Mqd8grrvcIV+9CXiAgplJJ9YKIjqwD8W+T8zd8pNR0fbFJM+COQylUHp0b+AaAbzNv
PsBMxpwirVcfAGF8VsEn2hWORTprmuMOSkWzzh0AEfYEIS15UQmviAGgK6oW1eFnQiCL6My2e+BW
gyMGRjQBnv8lMX4+eXd1tCZ6VK8BUTjub0eUGJX8yQRas/uCaWiu9CpUkbPp5SN9OChjxL6W26DR
l0ps56xhVYFhCyF7teXoXwyVEwqbh78OIkFT7k10YtTZHi+5Nkn/KjHRwle9EVNXGMILmtJQAF+m
yCXop5dZ3CqK64nVF30ecNgJGEfhUzUHHbqb/RCBkokhDKlY10DGGGVkmFG65d5QqYD4GYTTA/Qm
sVhVF8l8H+re0QTtkjKk2DQXnVzK0pX652mWU5XVfTAzR9nNOEqoEtHV87JZiPgN3ktnQ/O9uPks
6z9BtMj4LmOh3P5zyyBY9ddlq6/Ske56ltMCY2FtUXkPApWkwfLdFs3hEC3F15PVssQv9b6IY1iU
Q9SMrThsEbLEgRwG8os2EYC9mDa/os7jzbixFv7B7Es4DCkcBGLdJS4vNKFo8bjsc05WHI87P7Jv
vt+h908r2k4MMoF0Jdl6fOpWCwf7FJt78GNRaUcP7bxlrGRmvcyhgNloW+o/BfHtBMI5zy0NOJFs
zgUF9iMLzfe8j1YVTMTgGJ1zN+wLx4zYKxqCRzRdXDipAVSCA0AdkI6paMIqYm3GBA+Wj1gLNAnr
8+BPk8rbN28FEcgiSjqJCYJ8wWSylbOlCQ6qqjnN6BtNg7ZFwy+6KEJpNFQdACJSIRZir8tBBips
HFGRG7YCnbCpIR0yKSOLd3H5zGqTCBGnoNhjZVo+befrQcCvK+5lB+K/up8AJLM5nE9exoXGA21g
Od6s+brzwBPA25ojK5DAjsbwe/4NWUv1yBenz3EymDmTnpOEtdE6XiZkaxz9R3E/avb119LPBzj4
8tByJrjtXi9DPxhBFjO+ehL1tnqOTRj59b+R7vZh3Ygz/dsVsAH0ViRNsU+/ie1PPtPZR9YlYPJ3
R4dZNP9NHmkOZ4WIW93XOU7AXDFwqLc+F00Yuf+KINgYXl2R6EC6DlyQ/gpYpzLC2hLygJBFFvxy
0VvTqPTq3Hsb3cYv3/e6yg/9NWCmcIq0GrGTwRqNb19h7ZH2UgAd75O0SHMhYO2O1lvbRLZMiyQh
BBwFolIn7ABgLMHrw4r4QfFUDOUL4odIbsb/2AnHUoCLEp2XGQmkaKYynaO2A8SX3StJ1+aQqlaK
ENPvvaHc8fKWJYPNLgxKFmrkFt3ZNsENVc1GsS+sXuGIFnXSFSDmLjUiWagg1qvnHNND0tn46saI
DsnyTWy2nmnowgI076EaWfdR32dFbGC6I+HZkiDPaIWxkQ2J6mVcL/YHKZtnCStRgHRUdT01Iv6m
IRonOA5VF999mS3F9hlWhExh5qIFTkwNS58Gcy+u634ObDNd16etkIi29G4cXjw1g6jlnsM7cvFI
6MfwjfxFmtkKEdAVN1cRjz2jqiBsU1k7/EdcMMJsxFXKGbr6+KzBaGj1g51xUFOjbfClFbFMt2mh
i+GZE+7WQOAvEipJRSTVLVuNyXgyUoofTWlI9nMv+9spk9gDUxrtYrEwKjiLw1sx303zGifzEC/4
m8KRSUEybD6tIpfUlIh43th6pwwaqCRaIrSzBshVRHO+jqXugaKC3jJdVHOD8SFclZDSWCnC5wgA
pCgMx1o8JDdCYlYcORaP1YbF3hSD87sLjaxr27wHMlYdlr5WctSF4NdKbMLcu8W4wbZjT+Py0EMS
Ui7v4NIKrW+uAz3uL1gEDdrmrWUIBU+VKaPr6EzKua8G/L2uSDWRU1jQuERqa/gJXzgyr5i3IIim
moBNs66s8xawV6cexPY2ZsLDQxkcAaSZtoZLrMZaYoHvXVo64tTNCA+kO/Gj0DgvTVEDQkQCWTeF
3c4Vt3V222AG4PGLRhIja9lKV0CU8X77kxEFQZE2FM8KcRkTI9+aGN1/Swozv1cTVKE4TWmRbSRt
HFBemRyDfV6jUqwFsG1h8zzJzu4I2SojpfSIr0HAOg8kKfC4E+AaYaVLyCP22tg1vZuhgECPffPr
7M9GO9E9uVH7ZVgl1YGfdUsX3+rhRFRjzu/u/K8InailtLVljx2OHAS4Angdov5g1fvotSubhbxw
jMr2ijtgyWHRRoWkxJn9UU7DCgc6Na603pLR4vEgziF3WELuQV6nb01i9hK38QeJnY/H59t59PDS
o4ZPSM07l0iE9kruXpSBmgCru0eY68DxAI8jhSbjdaeq3f0IYtLTojOp+HhNImUIZGlkU+dLuHML
xMbmDXfwe/+vlA3AAfuRERHQX8g4P9Tf8mKYiSUpj5gZ+PVu4MExVnQZixq6eHrbnr4WZ1efm7B5
m+hpGV3Z6bq2hIWUvb4OagELSfWh5jPSH5urz+5+/Mrr/cA0dEleuThwcZR4MZsFQv87XSne98Gr
WZnZRZI5WyppU69LkWHpfSDQ92LKu1JvYtS7VAKRE6n9Ch1LG18FEvv5hnMcQkD1eazGmdXCqwyP
GfDLOm3yToBEQJXjVn5G2NZvp+bKsF19JvCanTnE7XCNeKVpD/qGtR4+Nk4PzWEt6I4spy5jmCws
3aKQbyLbZUIAjCZnCnHhAZRTUm2Wz0do8gop7JRLYqUIpfHVYkXwJrWpBZJsY0FvongD1W8Vwdnl
fh+8ljN7oGT60olmbELu72+FPzpxPs9Zm7kVsLGx3FaRrceKW2qtnyihHePKDYMMawcl8MPSMuzS
QsAvdoKoIwohxH1dH/HmmnFr2P+FHZdq0xWVQuc/3Oivbhl9G3FGAfYwu5u5LmLhYzLrA2HNK8Au
wCmZhwEiMs4Yv2FLTXSGqDHGjB7xFVkInL5DCAzHugnv/E/lnyxZKWwDEd2bS5GOt5cBCtsV5d4E
U+v7aJN22p91zFh6vwV29B6wdzyTgyFNBVqQk3vlZ2kL94G0rFjUczs2XbvJafz4PaGS827gAoiN
33wPLuer2szSY/kGabiECz4xfgyxi7n02cJkTSn3U64QGXKbVuY0+p2CdsbxDj9OA/1fl4jqEI0x
RSa+NEZ9NLyfZX+NLuhNmbBKemo1DCusiN8DxJtnqHCn1M2ssmMuXz7QBzgRtrr92AKfiQDqL9dI
J0w2dT9ZUClm+2zV5TnkmW/Jy9RtYda/2tw9kn8w0oCcXiT6Mo69tSXaHcRWnj39r55sgS/ohbJ5
4yD/3Zooh6PY/g8+IF6hF32rOuhwBfnsG/eEi5XY/3PauJobzC0wcNS0lXAVDd1HhBnHaxXSdV97
VBTz9KjuImWRJ8TR5T+cEIFt//I8KC3/UzNvVhDzo93ZKubvvMeaBe8DmP4aT8RZIJ9w5eGaqfXT
3iJ0JVoF4kckz3XsCIF7SFBuZAnHclrzmrlaArSlRaSJzjE6r0q68Wv58VIChuLbPoPUOLhEC5JR
onAmtM+OxIE93i0UPjSh0h4swj41dpI/zUpFagHxGHzOJCmI3naO6+i/zeSd+j/1nkY4+iFSCeSl
qVu42eF/5d3HF6sXIV6XzraZrhN1dpti3jgoZ8Aess59G5HaLeOHT4TjL53eLk7UurBdGOLxYNL8
Rgpv60P4N0RnWr4fqGG5nlfSs2QLH2QFdz5hH0WRT/TeC4FlcXW6/94q/sm1Tj+1JL1YEc1V9zxj
u3JxEWWF8KdkKZxeLBOqLoSRS/nAB9RTT5YYURubZS0KMp5F3e8jaXIWjPUdqWgBUdcNMIOEy5qW
a5Ose+NANYfv12K3z95Qzh9z/ukHzDu+ptP0qdaOvRCGQu3ZgXNX7J1WBGJuL0u29RQ8zb3qC8yg
pI1rwX8VPrh3O8W5FlgUloRsxC9RkR4xr7wQGAXVw7f0fqUZsnsOJXkmab+btqSpDmLUebC4ztUW
IIhN5qXSOATXZCRYkqJ38p+v3kSgw63R41wf5YRppHd3QO86MqMW2vfJAxhcmJr06aIAWqKTUbG5
wfGnjBAoSicw16cYXJEdnNeF4KkH/K6Koi3F3FVUc55yHIwF68aiLEU/8QuZXc2Wi2DPYQqw7pxT
vjTmz/+2/A6uW0oO2/YwOlvdRt46hriWbV9ZJiXo5r5HQIgzgZ074mgOIPL9p3IVgCD8Ejll5Kcv
V4kMW/mWKeyZQ6QQH+L+w/6Nh4XkzoxBhFPb1fYBCltSCXxxNPU6oYGSIWbS3uxdfmuXvugY/x+B
WPRVvnK6R3UDn83r6cDuNVbdxEFwiPIvJYIqZ6mYytXQktQOw/ITgCnMmEOjymb6la2GuiGRX3kH
YQSbSee5IrUEIpZ8PeoTxHPPJE49bh8J9HgvTVkyxnzdma0h+CuMJSeDfH3A/88PqgwF4JeDrfUG
Ett5RZVv9XYYO4bjjolLP3dQXOZG/7UW7Xrje9+xCkXLlpcjfB7ntSWFxE8B+eTQPzR9UbTBV+k8
QcSGGZEXsMoVgHyX/E5Q20P29pdTb4MAPwIt8/iCqvzdcbzYZH0sLfSX6LCClsNZf66vZPU82giO
7S3XNCLgsnMmTiJqfTHeB3P19TX3/JEUfrjRv4QpjKEhn2eg+N2n18wv1vmhQEw7SuDZS+6V+0zP
zfrGDU42OafISlZDQQRuwu+v1TSPbJucZ2UpM8NOlRGSog/6Z6UGJYeo6bCrLxdETuWFyH6COaz5
T3jQFhjLEhW6XqKtd37yc2NHYag86Bc4k+d9Da6/CaOf1BtXIl9JYYbefsKN60r9q67gTWbWS/rB
IVHzrp5nYU5m0z0X6pIiUE2EiHjWLcsKyjbf0rIQbHaTXZ573xz/WVxqS0vkJQjkuEVRAZxYgT+4
SyCZCIMWfBYgz2tueQrQ6carg9NRiPArHrw997aYmatgG+Y9TsNO4yoft6DsbayTsbom+6Jc4mms
AgG4JpXhG9Trbos3qh+k0c+3nC8AnlEjOc0Mq3x6oCSTMTY+usryosJmspPeqt9tbA9TMMPD12tM
qtZwUABx4WG/tEhjW+iwppCe4Ts27zFxTD0DzVRFN6GBrGEEDmP8FeAW9EQ/zMCIJ+tlewJFpXao
COQsg2Fsy4qBXu5nkwExhh+wksuzy/m/cGOnNab4jxMRZ41LZztMx4iepOmm1AZuDyUZVh/FzSzH
jyWjZ1QhCOJ7fRD20pdMAf9e4ygdiOLwDhFMSwhpHTA4hKbU+78Uu/X9sVtz6+PxUK8YRd5EhdPg
wdWe/YdvbIYC7kFTrXXly9wJ41OVo1bkbgf0+u2mwKo5w/iWJDWS63BxogktWTlALM0FlTkKuCTH
yzW9McibZcCNCzVUGqAQS6aY4UsWTLoP4ZKYa+r5ZtBdjvkfJzQzObgpOnyv9EatUjqbudMCaX4+
esVGIrttKdw2xTljXvV4jyYIMPsYAHj4VIE5F4HkccMO+GDlgmcHA8LvZSPWzeSGx4uctVXNtAY5
uUnq0G6hcm7S4PGyg1Xyy6VVIylcjsJdwmF3mdhCFWw44Yv0yYAjeAkW8dWMMNomylxi464f0Bni
Bmh8oX+9sZQ4DEOQnX/X8k0V9MPmpXYOc6D9JEIl8qZ8XyxdoC4h+Kj/KNJETYCD8ks+i4OMDnGA
gnJH7DR5p6duYrOVtVqvabyetT6RNtp74h003Gx/N0qUAJDew3ZNOh0YfAI/yoeKN4ixyQIuDYFY
psqEfudx5+xzfshmW37JShJJry1pCZkjO/voaWggd/GNH8wPwzaFfzB70ZvG1DN0GK4r9gpwi+fD
8VYqlvXNvwByDzG61Y//Wqux9tMfVaKF3rW0zGmGQdR5pMwgdTDa3GtECm/BWZ57yiHlwyyHOk+1
3LpY/KAx2k0XJ+nOTCw2X+KSLw6YPjKdyKWDHPA4iXkSbFnEumyzy2FQp1MiqPdev35AGysTEB+i
Bg6cMlsrSziVSiUA8aXPlPjvqXcZ5u4R1ysk2vc2mk33ouqvKBuCLdDEUNCtzWMS3V7dBKmCgXrp
tIxKF2yZF8Pgs7rs3wyzjYD+l89qFFmZbKS+QRiRJ9+rc5KPWaUFKa3dwbttyhrLfVAjVCbvq8MI
oCSm2DeZD4mInyf442nTA39Gn4J3x/RG4FVpxlgJk/DnpOePmLFRjxKkYZCezC6MHgaVfHHm5XNl
YURz5rhNg7L8YTVHF9/VS7Shhki08jDNZcigAywOjEd4T9RqX1PxdGjjZbGQRRoh02sZ+YdmPDd/
btpDoUAtaP18lzq7IGmlamXqq5fjVnNZPCq/rcT7E5dAJhxoGVSDzb8NTfKGF0Sw/UP22IoBgP2k
zTSOOujTZGxe+oun8OJ1jhuui7jwflMu+4Z7fJ/CIRPoPtrR0baDtWikm0dHGwTV7P9+iEWlqgd2
zRjjLURBflI23BW6QqM9Wds6k7h1hnrPGgHHvH316L3oCcLuV4Cfonj2wWS/JLm+gS2fJxJqc8Hx
+N6fgNeovm/+jt4Y6ftaGLRSComsHVNqBtqdYProci2Oy+BmdlP0X6L75Q1O0ciV5Q5C/dTMOY8N
sp5Pwk6dkXE2JA0nCf4zm3aXGYclSZJ0pBvY4KQ1xAKFYMyMC9LORSCOJPZ0SAEswtBzG8rOfblw
u6c8jDpyZyuHQoMuCGfqSwdI383IsH1JB5NxZQ/TKZZduhmMqZdXcQ6ZgCXxm+N6n4HMPdVfo8lZ
J14BW55XBjUzAFpxj5aG0Jw/a6VkYvRjkv7xTKLz29daO1o9nfaJwKRSxmWKdXf8hrDBuKiapawe
jZpR9nHq6gBZSFMw6Ye5dQrH7/Jts6H3QcdyVdHJ3e3XhGdwyDj9IrFl/dKQX/avp9EMQCfHsxDd
Je/WeVKi4abZUUki6gWg8YusVdL895+ntqhMOMy1qvTtg2YlN0zUFPZxf4qaHyZii7/yLoYd1YHN
jLLDaPsmnVSUyJ7lle4psMhJb6d9lfIXM4XTHLHSCJtkqIHbIVw/mX46cZxsg3RYNFzBOMPEOfQ2
tTZA/Qk0CvBTN1uizD63KNCq4N3+jnsp9s8o0cbkXGt+EO7TRS8k5or3u2bxu8nGRCvFqKcUIlWJ
TbIq8YqEl23M1fT5OCG7uDRtGSD8xDxCRzTdfZ5zzBjcc6VXR0BaQPoIsqu0PMfSCwfK8x6ztZwb
7nspb9/1Z/bXivd3jCQxZiBptpcIbQ+wDsyiFQBGN6EZ+9PTsT+zZQ/xmh9tHdMuV1lAVRINLRMl
W+G3/lMt31EJi/9vvtvPdqKQ4HfppKo1EOEks331nt/C7ig+ZWVzeKItNYfxhrItuxycw2Uu8pnj
hGL/jMaYUghZVoF4aSazfCKvVUAV65tAWCxdfaU02koz7ISOncKJijo+R6SCeY2KaLq9m3LiNiRe
jn8DZw6f+MjH0W40vKJm543ROlM19M1BJs17MAbTowHUNpPG8VzQoZlklVkPCB4/MhUfVzCstd1n
wH26/UwivM+hGFgAxQ0NVcmjVZ0A4I7sXnHz68sX3pYWZ6WetZo1Ym5oVfs190EeFgDnhM8Qie2l
MdMIr67exmfFtH4reA33TlZNfMxZ2zYSYPFocd4sUSKzw+yUfSqUrFqfMmS88o8/yb2hGKy0EhIO
5OyhHZ5wz4NpZc1IyrZmPibB95ZbGAvS48jXQEGXqpbPJkJZZVG6CeAAlIIon04OLTefdGWxw8kZ
qChRp74w/6JPMEncD8tQlsg7IAkGfMwjUzavce4sOmYHx457ZBQZFE+YfT2IDtrgS+5WD2Nz2BJ6
+lBsw+Ni7fZqVLAxtstOuZ1txd7G2RJtQIdTD4ODSrJbY48ieA8TpUsHdKJrRvjw9V/d4qZpKmDS
2mCsZGOoEgVNG32tnZSkJtcRw1MCMBrBesZnhqf3hD4rKnyVCEp/Rt1aiyWqxIbp37rxjSkJeKzs
b1MjjVbdKchrbcXHoDqUhi/ZPs4thZoSVwK9lpP3qtry4x4jBVK02r2FkBwXXyED4JCG/OhD07Hk
m4zMZafOYaRc85QmwIx+q1d4ZXkAmkNYdQacf6mSog8vOIqTXPw/J6LbATLZNWDO3gJ9RxVr4JH4
/BsxKWR+Os7LdUKpTnhbl0oayV5IvqZDaqgDFOeu6mZdOb0K411GS+uhP0E1vlQTvhF0aOTI3zm2
KOUtIBrPPZ2EzxQ9Sa6C9yFdMH6mS1DK0Nq3lQSAUYkTtnI5IY3h34R2k+hLVLOKh8J3e/jG9JAf
bDJuTTCFkb8sR/h2rfB9ISOXInw0EtAtxfw1ienTzCIqmnYDFyIodM+/kSjotq0lANVyvyI2k2x/
T1o9tN2XSYsrXEF59YmuIjdJmTpPeMqDuk29Hpsyo56nqBthBNZp7PB4dz/LEXw1NgzO3mnIgQ0Q
pdDZNYRDjZYOg1h7pBWdQQUgMYtSsTP0InGQ+IoiAB8kyH06izlS3JjenMP3OnRqu+Hgf4+8HUNy
TOo5gx0544wWE8rfWaHOe/Kr9q76WO5l0Xsso+j8RHGXuLOygDQPrjVQUs5wOUrBYsoqKOKVq4Dr
AVm/QusnYa4E7j5Fv7ed0AkP825+G83zibvXh1EZzFcok3q3DoS3LG8cSmxT7ESNcTrPNZN9r/J4
CSqULdApXYHiWY23sn5hwr1P8eImxanfW1yd16Ghl7sn1J4PJoKvs+M7ALK0lETZYHiNM/MzBKar
KUc4j1/yY+bwfxLZufPh84UEg5jcYF+fZBvRhLjmhqrUB1xt/51wGSyI2TLMCZ1DXB3aGYvr6uVU
VwhQyrF2iOHFtLPn+BnJD1vXk+Z87W9u4zFisz6y2P7H4AcOkjZE8lllKNlUJD1y/L270AIWfKs4
G2+KawyEIUcsHSAcFM+iDAF9EPaLG95wyTeKl7jwdBDkJZruFDOF2LMth+zbuDV47Tg1iiXIrXRY
Y9PFrGs9a8vZF9gLZhBtAR1OCjHQMlcCCt6g14nLJnrIzPscjzSfHdH+PhXTaiVkSAVzROYESf46
S/7HktN7fOYWjMtuheXJfquP48xmu7HfJFCyPptwzJCmwjMW/9ovwwcUafnsCqhGv/FKZf3o3DiP
BysfeR/zzsIoCCsUNSVLL/AKvIAFGEon48+IKavPIrzns6Vj43fqcO2Xz6UZT1TZ5Bd8xKHlJb6U
lV4bvE7LWfAff5gvIn0Rypts7NXhOil7PUxt6kPxKLRIaRoarB0+eB98WDcD55PUmMzzstWCP1ky
B3mEunzxY29/0154OC0EJaTINzgOLcKxjACQYGLPXUaP+HKgRm8zuWwujlJIyTRbmKDc7OFJIQ6J
fNtfUAibwefdhLP6t3af2+xjroiQJcfLKapkVFhWQRWSAR9lThd3HyYALNPR3K/o/sN/YO0E9Hho
3ruDyHfG1h6Hbq22wp7B1eVeqsDl/RN/EqbWcKlAgWZqZuM3lw0QAOoVlM+J8+d2UYanGqt+GDrr
xWgFPHsOm8ORbiQfxxIUuiFvOHqP8nfRoIc1l+KsPp5dIroZ4FKR3givd5i1AjMco7llpYAvQbn6
VZTnQyJHNmTnvqXN4dHGIiuonwJb+TUQKVjt+IumxJ8+ng+IDEnoBmiKxHte3AdQDicWoPNHTUcp
maAxs/VKM5oSrouqC9l0M4GDZa8mlGZik+cyfWPR60CfgnkIi31S1bBQ+lbISpb9Pek3uXb5Cdhm
IB6N+yWhbrBFmHAH5jJutxLd6SpEqLZBoAB4/BezTTiWJMzBzcCDfTHHndr16L9p7fX3tmaw6ZeQ
b0zUR6GdLDB4tY0VAIUYKuXWinKbdI0OG9L2qwFLmyFF56uAKxkWWriKKIYcrD6RKVsLU+QK6r+j
9S4EUgi2qSRxaFcQku+5R8M3mvWLAnaPrixHms8AuEwgZZH8FD+DLvBtM0b+3tW89Tee8PjIPIvK
6HLAKCURloRxHegXZl1ljxMnGD2FFoUl0SkMM2qNfjotTtLpgr9Bv26skuJan0agDRlv/i76Y8A2
81Oh8+DSQpTrr4hoju6FfLh6lWkBYUPWswj2Fucx6akr3ZwHPfWhEBJ80Nbdv5CmQEZTPPsY+8CN
uFw3+cFVmnzzjmvGFIAFXDufbu1JKcwh4T7OV1rHB/HSgQ0VZqJZjNwBtRrS82MCoh7sDy6Ta/xd
QOiF2f+sSrdwc1veOdyfw696KNVoDo96V9g0rfbMpIo2JDsOVCQPGR0PjYEcJTJMG14qRx5UwvS8
+oIQgItdNMtrZmgOE6MWh2aWznxYJTdXEOLsoZbtPDpCHswhIMaOFmf/fZ+pwgNa0oU+9Nly7Pw7
4NSahmygt/YSy4/JQqQHKexMCTv/X7bUPq7vPwC8Wym3JP+TB7E4AFm9/FOR4qHYM2N6Fu/sbwUU
t8fQ3Kzyoy7gzeExPZkKMB4mIN2yoUPSSnzcpzTSDvejx+Ss8rBPNg1ckOsj0F0tbWhGO/dbVGYW
GMY1RHfryUCZM6sNLHDFEuWERLvbjZ4QkxLwK6JoEqpxxs5qNOrYRiQ9DaVmkBB9VnrIqC7L9sck
fKv0AcpcBgKBlwYsDBRHAjUPKvVMFH7gIYeepSMiu5AND1anK1saazYsZXaTscZ0OxPg70YWmDcA
0KCHrl5/lsllJvxkM/lksd1dUBXE2ref5Hs2/3svSulzkq6Nf1WGiydGQxvsOkLhjj/Gbm3xWqud
vI0dZA3TG6wsS7wQFlNq6+wLZBaGO9WWG2q5P8b+/wYfbv0TBfq6BAA1NTvg5JanixmkqFVPQ9Pv
eXgdlE4W0rrUnCJWyW8llhqRP8qydAG+BXyn2ES3CqvOFf9cjx7CXgb+wknEeiOJY7Q6kfPXzIl2
wRHmZNth7TJVHg68EXyxUELKdY8fnJtA74f9lv5iJgw5zdUk1zDCMmIBhpKWnDBbGQjDaE8fyfpn
zhQ7TE+0yanaOXixz0FT0P6aqZZWzulnHr/DVh4Xg2h18NiQTMxr9T/xBxRVxi1mOf4o567P/jAK
uMOjeY+v1R7lcB5Kh/Aek6Vi2ERB0hAwZLwysg5M2kMhYjLjjE8IJQahaSC1yTeWBX3SK9gYWxD8
FuHYFGkD3v2YrOb2aB2i5sG8ICDmsBRSHASx+AGTLqoWG/ALssYlAV/QlBEix52+wkZgkAGLVb6c
pxziXsPgmhQNLiy3NDA590dRbWuzJ3Bs+r3eNtB3Qz2ijKLbFOq8pP9CFCVZVf4Uo0/lm2Oflal9
w8czgWHgpHIzIudWyQwaw9smBmzedlymnylLswsdokVIuoaoY2nUibIsixG2ylXSpRJP+xPWadha
s3S5B4QBUzC0mNT5KQx7nZyRry4k+P7zsQ6P+vpzxttEfR1zIgEeKFSRX2plyGazrcreVYCGKgyW
8mn7cHH0nRU5x5sd/GGF95hLD8198u/PkJbWNtJd9rfkHL5tI2pjVPHKBs2WUVTIJzqQEqv+nHv3
hOmLFGOV+Opc63jpjQzSv+Z5l1JaQ+lPvGgYcCueBcxm6GKa/+E8GAsHqdEf/SdJXkIzxJz9JzN5
mzWvc8g2o58Px8FsjSsjpm43kixopECoMo+xWIkAqK+GtofEY3mt4RuCkdjO1MQT2yuGTcG+aPYH
fXbr3i+fqWIBzQHkYrZeCI2kYN3Iwg6dD/6KhHm+xma0BKDVstyruo+n1Fe1rzpLN9kEQc3zklk5
ybym/qEGJxqIjhjHNt5a4QDMsc6AYYDDfHMqczo01OrrAKFQo967qP+/1BoMqqcRpwasSnGPDX6T
XIhFahiVNHGX5bHGZF3DeLXI4DabLcIDQbsH16MQqqp+hRWo1A13hpwzC4TV3F1HgYEFEAtvtrsW
zinIWK4JvGhM/xKiaO+CndYNV0bEX9MiODXEmQmgqzhZ7YjhuHdqUfztCTT1+n3ANavijweLYflZ
4+SwNqEdoca14No/cLzJbwmQvlOlvowkOQtsyLCtY5W8bo46Y415MWR0A0DjPqTXYKDnWeugPbP7
jrfR9ohxHX+z7hiHuXMDiaOr0Q9gjMXf/Ow15Msikk6574V3owgcnnagpdL7pM8jVHorNXDBWZ7u
Ime/QgfXip0tz4iNJED8H+lRimZBMikXeafxfVxQjze6962Sdc2FlkhiTM1rpGVhfDyi19JdnCvz
Ukb3FNprTCQrpeuiE5+E+/q1GVlgGo4N+LakMKnY8Cgd/U28PmoyUp+wuxWG4t03ld47sEuKSSfI
8cU3mke03SId+jUOAg2xWY+ldXtUJPvbRV++Ewb8jHpDPQPJ+X+bnXZTPQ9+SBNiSvuWOgBqUTqT
lQvdqI+evI5LtASgsfPTC16dObos8liNIuwpJwmC5reEd+95zZnhkrXRJmM6a1Q8SdacqR2AqKbB
xkorS+UOtA/M4yNZ3J6BohT4puuGrxN71vaJyB5/ZpegxFgJYtHjtIKuHFvR8s8Q5tO9NFZyIbfv
bD9kOPMY6SJSqUPEajZBc0oF3n0dDDEhKchRtXCXvkv8QpTm8uAn3wB2HRHxHNfu2geLyPsznVbi
dwEUBiqFHSDVi6d8f7WRXM2WsTtcAKQvLdG+oEJf+PmrnABEEesAxFxNO2cHO0HrFh5GSB9/Cx0s
oSYd/ZPocIJfbjV/baTAGkxH42Esy010Hj3kUgIQmPE7EZEv9VWjUy+632XHhTJHHGXxVKq4lmn6
QJwa5w8dPe2Xy6fbtegif67jKFW9cWnqLG0kDbtWwButsE/SDddf6twQNtxe4i9bkGuY0g0XQXye
ELjBhkhJIiFAGq8LN8jjtLcft5z+K1YQPnnJOAL2WwmjhYi3ZRC1VGZctMLRQRbU379/AF3+RBXO
COKvI+hGEiqu0m430wNMTzVcZ2JMT12cWcrC3JaCZhAr4i4LhUEhvo4wPbLY/ecOYmAhAQx6jo9A
CrSbmSLmg8QPnqMt3+EQyH/SQCdr+HkHjE44dGqoH/5Ni+IJkmCfc4CwerTVyMiMU1JGiJszYGEz
MKp3qrZu616xmCDyImZbzWinYnYVr9QAHNLwntwa04DFVmJNwxNOfY5eQZVAtJjUkxDHMxFXJu8t
02va1nsNoNQ5b6awZYxCNqkanuDEDlw4YoDdxQSxRH6kriO1/62461NST/TbGP9n58or9kjZUNzX
sL/xk2r4rNIuYiTgjy7THNupuxq/jf5hfO4xqBMIoayCH6pmJcTP1ra7SNsZ3wZvQBmr
`pragma protect end_protected
