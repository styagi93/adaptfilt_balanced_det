��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|��VED�׊���nK��h��tI$�uuC��Ah#�H����"�q��{�E1�O`�*w���f�ʘ!E�����)s�'t]��55.&9��̫tn�SL(\�#
�k��jIeKnD��������U���[N=3oB��$���I��J˃�'^�����B��� y7���1&`����n��"��zT�֋���s����e�B�H(|6+�L�O�[8	��F�~=U�k��C?u�ep�,�o����4%_SU��q�왡��z'����u�*4ՈQt�"�p�^K��/���N]��'�k�ȑ䪑���7�Z0�}I���$3�y��^���T����wu�Ts�xp���%�h�^\���m����<����÷<��'q^q\��s)��P7FU�}��o�(=�j�w%�I[���+�J�mr���@�L
�b~)XR�I�� w8�mz�0tt��\d�Y��F�/��q�͋eN��?��T��Qu�$+�m�e���&���z��Kʛ���U�+��@:������lmCbݦo=@b'�!�hF -�lC�	�tn���3[��<n�3�;���">�������B�]��8 熎����4{���Y��%
e/�_��[U*�J-���k���++#�o�Ӏ���� @�U� K�`wNl�cL�qEk���YfN�G������#L�K�L�&\�Y����7��-�y�W�a���C;K�&N���EK���G��w{p�"sX�]����ʂ�H�}��2� ] {z'y�*�c�ӛ�f-� m��f����3	0�앿BHlVP�?��f�A�EC����bh��Q��+�s�����"�xR���.3���{L@#lXf���@�~�/CZ&�@}�Qt��<�i�3��
��#lC������
8GS�����5�D{n9��=�Ll��� 0)*����TG/���T���	�zG2�G9ƙHax��20�X�"Gh��~t[���)mo��%�6Yu��0;��5��W�n[�dB��r�+P�J�haLϓP�35��G��� �`��4E���+���J��a:J�t8��i���.4�b8�n�U�	�����l(P��W��p��u�rGM��r�ڷ�U��w|>��Wj��jߴ��I:.���il�1�^d�X#zHuB#I%�?.��N�~0�V�b)Wyc�z�)K��ǿ$n.^�.F��"����m�o�Q��@1IL	��,�+���A�C��Q��{�s�ݓ8�v;����,ׂ!̵>�Y��D�J��1_z��r]��Ոd�-�э"��[����5��צw�z��D��M���$�=�`�u�|R�k��V[+�G�%F����k	)�Bj
�����(��f9,���������;
�qf���G.�oɣ���/�teo���ޟ7����>��(���l^!���]��_t+:~��P&�HdN�:�!��o��v��)���FP��̼c��?�0~�䬧_�#o!�V,B��i��V