��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ���^\d��l��m������� �P;N��I^Cg�U�j��3g�o�����;P�П.�����}� ���T�[�͡9}�5��M��AY�?�����4`�@�O��Դ�"��VЊz�Y��O�%`��S���s�������C�7W�kZ�?}���g�F.1��s�}h#��?<�Lㄗ#~g%UA�gI�;��<ص�o3{j�R�t	��į�
BȆąV�D�}	ό�����F��ތ1��[x&�#��!1��O�R�2���������m��W~�T��S-g�Ⓨ^W��質h����+m�����Jñ��1B��mx��1����s=њy2]]�?�� ��aGP��:xc����A���b~$jӄ[+�}H���閕��Rל휭����A=i�BI��j��5f�$��V��`pr!*Ft��I;�I��'v�@d5Ygu�{�O]m�۩έ��{�ͻj�s��)e��$��z�������yI�AX��إ�c����֞>9�>[��tB�� �4&��8_�;�y����j�o��g+�T�/�r;]�\�=��I�a���q±�d�N�Ĕn4<[�r/{+���z��V�P�͂=(�Ɖ �_E�>G}Y�H*32Р=��αM:͒�O�>�3��h>���\x����h�3�c�
כ�6��ν��=aQ�����)�S�
3x���*�r���1J�_=7n��C�g�9�>��q����dݦ)$ ��lWsl> .���>�ړ�^]_Bc�M�ᐊ ���������/2S-���EC6K���u6<�In�%�f���{�s�R�Z�R��vb�6^$�И�j���YV�M�`d��C�l��g�2���yjb�må����<6a=A���G��B�̱om�
f�s�Tى+�F�i.X���;���5���P[=�P�a�U�^�lݙ`��d��yӃ��ƍ������j�z�1[��+�|1��I�E�����
᧙��L�����Z�VK��0�� �|^�U]ee4T��):����L�}�[��*�n��,�&qb%6�*N�$��v��R���HH��a��Fm*�Ģ��z 
>�j��Ѭ)�D�{M���������w���R�B)7�]G���L���5H�n3��$��Y8P�X�5�K��W�v����a*-+ �F���'�f7��Τ�Vf���\xqais���]>���b�@aa$���8�!D��f��U����,��1��[�U��a@6.�Y�+�:�����BB(�4�@T����׹���/ҕ��Q9%|;��.�2d��5o4!oM�`�C�o@���&YM|$jR����,fƜ��u��xeib�m��D|+�z�'�;}�"Q�폭7[�؋bp���=؆�_�)ɵ���%9�1C����2e��Üc ��c@��
y��:S~B�����N T�J��y$ֶ����2c��\��L���
�������>��C�Dk�7%Ǚ� c0���k8��J�4�V�[�A�?�:E���iC޽��%��Ik�n�R�TwU��c~N����=��W���'�/�j@03��p@$�%1Ī�'���]DQ��jf!����W3
�I2!���mB�R���t�y���'�����i������X1x���{7G�Ba� �w
ggǮj霕�ek���Oy�^�I�/�^�b������;�m�>�L�Y�y���$���k;N��2hC�S��M�۽�ר,�w�e��CV|�:S[��U�r	5O5Kybikp���;o�"ռ�-�ўt�sF�/j�R[�ٛL�D��5��{-8zb��^�+H8����U����P_��F^�A7}F'�|���&�cЪ�a�������z65�x��o6u�a��U�	=�0fk�Ͼe�3>\$�.�R��.)��������F2�E�2O	i��,�h-��FU�_�H5�cWs cw,XsN�+}��v�n�)K^v.P�����@]Ò��QjA���@�����z���շ����8ќ��ּW�u��x�D��D�e