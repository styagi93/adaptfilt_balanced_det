��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[���������,HP�E�E�^ޝ����?	�$���Yd���C*%��7���+�G����Z�騸�Ӗ~Hz�l��;`�9䠰n���R�����n�W��݆�U��X쯍�݈�ƕ�Zm�ﾪj��b1����.�%T5I�1�C����q[�J�;�n��5�3u]�JO-�s��㶰m ��pڃ��N�=e����L)5vr�$��3��Q��6���\H;�[	J�S�d�<�86U�m2�q`2"�r��y�񇪑���GTO��t��6Q �� H���>E��� =kuī7
��.�\M?"�|y�P^9k9����R���F��\��)�AJ��O�VJ��4��/g/s@y�{[v�:n�QaLޮ5�Ԋ!�dOgW <���
��CE��3�y���7E
;���q�K����-;���͖E&Hegt�J�����"K\x|,[�O�B*F�+��������h�74�<C{�;��6����y	��q�y�9�Nú��r\Ko���(5��E�3G;����(f��Ճ�.����e�V5�Ejjը�����""$��-�"�p7�|܊0&Ӓ�U�b����sp�LH�:w�|Y�2��{E��R�>O̫����G���ܷ%����rB��IG%�!NG.@��MU�[ȼ��I\�GΛ��v�Z��[���o�8Th3�drr��P:�Q�E���xv���JPT7cr�0�fwK xA��.�$��=�K�=o�47�x���<0�GǗ,k��1mc�e�}�%��4N�G���mK�0x[��9��X2.SĞ�Ӹ���n�O0��Kh��X����;�˼ɐ�w뷷y� �K� f-�����eN'�������gu�e���C����:qǙ&|�<H�������Xuž��u#8%4�Q*��}���,1�[�,���Uz>��y�4��r����8h�	����ə��
�
�����w�H�<�[�V�E�a��=.4v��8��[C48v�t{n���}��'�������4���������(a��bO����=��%��Y��X?T�uڝ����D�R�>��i�7��)R装hCI~���	U�~�vLPp�e�