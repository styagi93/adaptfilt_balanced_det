// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
zJpjmxU1x4bukkKiblSHbI8mkwAtcOEbOPM27mLqQQxB71z40CEU6ul71/Fp5FZsQEmagrxTEj7r
31qW1FdOtWp97Xw3we67THCQWF99sUatM+ahT8FT9rH002bkSuuv9KyRl561E94nRDFCqPqCXPU9
hnPro4r1kwgD8CemxoCYgdsz/UOSInhnPRDqPcRBJxZ02ZlekATTmXFQOS98ktjAdPM+N/9m1dTj
WHnnE9ODsoJTsqV8XE4550CTC/NxVZquP/Qq3AcOhDy1IN6fIR34xYWxL44+zAlZEz/t5+gLt0yw
hd5x5Kx5iHNtl7hcgEca++TZrxFVvIycKhw7fA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17280)
L70ztotsR0QwB03tMSfdP6pvasoCOfo4lIndCpsDOFUWWTyb1FQ5oFRsdS+/SFippbHA+/6ctqAZ
lEYclqi7GjBOeB0dy+JHgTgr5peSzzX67TuC31Ie4AfJZ4gcPQGV3YO1AQRKXnGZXWPY1/fgXVx8
FwkTEuNy4tu7kym3W3hG3Avdw4cGKorouVHqrSAEdzfMVOAdiSJmEAsmmXl9GI2r2WM8TsW5Fzfw
jyukii5aqYGo3vEO9wg2eSzEh4M9hvDImNr8Sd3w1APJ0qE+NBOqT0v3fWv8p5rTv1kavOeIh70G
ZQFcs1TG6CcPtEOnnGkDDXF0WE46j6LvU8ZSwU1/0dtQ2TEbjqLBOmEV5VAgvyF16DZlyX6wkYM2
abmNQF1hrNjW72Qd60gNVxWybF6CnwcXm/jncCRsF7sv8lTwk28YgFLKlXRsYghiTwuIgn04hREI
i9JcduCjpHYCV2bY1GBNEu+oA/8vrjRIZWqN9VRHnHLCVlxLioOsvrLiHm5GooOOreL0noEO0nbh
5TiVliWQ1ZI7qH2A8nT+zono5JZL1sMK/PZ0p2D9eOHh6en9ft0VX8+80TvupJqzN1Dq2tUZHmYd
/ebQfA+OvU5+F/gzZfIBeRYifra0BJ/Tju3FS3SJ8r3znglOOgnb2DK/UH78/HEg0M8Wdwn6xsBC
mCyzOuNy6u/6dO2hGY9OyBRp9l7Bu2D2F2pcTd4iHFKusgx/gkTusoZlO21ukrj21DV/U9fLCg0G
gwGAoL8NK4Gm/f8T2yebd+GP5IIcYtQgpc9vLVntU80LbP8fvkSlG5Wftyd5w66xrFdY3JMVoMqo
ol8ldd9v9c+lTshgHrs3fMOaLQETdvNOHoy8YEyA7n0JfzICdk9JG+tN+6S31pLJD/3ibii1XDjq
yq9ecRFsquQ7zHWW85e+KLSyd5xUNy9ZJQhxscM65vo4qM/3iQDLMinjiG1828a7iHhPA35r23DK
80mOQSDTq8IgoRYZwl2j8eu5KM7jo9z1sQOUx/+2+b+pczPeAn8h2rGXn2TmeWjrj4LCVctdVEok
ikr7UFKVAyqLQ76XDEY1ODfuKkudVCNrzwmtyxaBFsamto/6C0unLpS6QaoZr8d+pMbxQ8jzqvlu
yGDJWHvAQW9xmcqV0nN5ihE1i5QwLLd3sLcvbRKKuf2MIIQJ/qDN6QAf1B3WWBvreWFIN2bEeZxu
KbhdibWeMj/513xhALNEMBVYR+tZvBOrgn/U9zble+r2Yba7duBcFMczxcmQgp5DtuoxhDzEejZa
BzEJKDRKUXTNxJaeUodcgDJns9fcpFZrXifL1PQNAEeDfxyHxc8OxqJSebqWEIY75chgq8B1qg36
LLJbrF5GVJaocImABb7mw0zlgk3C5wqozPD291pLjq3R/YJSvwE8YNze7QYuqbsv1BEO4pNEWysg
van1u3EcGdN+TngHjgMySxxRbBFmp8waonhRB7EfDeDfDIGz7GDtqgF8jv5Qg2c0ngn3SP0QWH9f
+Z3XSTimZmCbhSSxO2JCtaU4fMIzowzNHGNJnIP5SfWYMwsyewvQd9OhfBuDgDVqUswFKmOGY7B2
squ+aBZ5ohIBwU2eKx0Se1N/Myj+9Q+m2eQ8WTYtpm/5ewUsHqgCd9TGcvuP8gP8QPRkd2gIlmaC
F8wJtq78pl5QtTt7RoupH6tTQSJsl8U0oRv4xrfa59JnZq/ZfrF1rP+Df4pz2xoO8/4OEMkBkqeA
P98n8eDNmUEtyOkA+CZQ64U09bjTZ2fjjUtlUDop+jo0lFzjhXS1A68oYOQZrXLNsAW452p7sRH8
5UJ/RpacEq8bKGd0qcLlhVAsgAkKl/0kZk7a1E3uySiJm9izAbJLj7clZJVeLmXJ3G3kXPTkQZLd
9lJ5RohUSqW2CMsD5LxyifF79Ao51XlHq4aRFu5RkyNg0hTOoM2IRN2KvfZ9k/QHlNfBPJ8RiWi/
hObHFIKQJH6/eV7EJIqwzrbOOSh6fxq/Wqsl1HiUyWPNdQKmY9vabCOba80GMn0bcALzjaHKCkJY
4aRaDeMX4abZzP1j081hHP7du1pKY3HOas/ApW7Hn8KO9QpZkCVmVji6bIERgPSFejA2IE+/+7cn
HbObCR0jkSoxon9chCjZGDCEXXzRD4O89RTtpNxUwWCr0LYwPdSQEEaoLV09o11Motibt/ZJ3syO
81hmc03/YBAog9DYltRUkk+19ie0WD2GgKHP5MXbwVhMkATg6jSE87zbJ69h8vVHsEggxaDdr/q2
zzA2JZxW0jorGhdMd18NQuCTf1cJA0TbxMFYFUKBdvhHvg6j3zyRTtuA5BLxa2saKUzGlvBPEXT+
BGkSaTLhxOvCA+oH9XL/dLF4uAs++xd+aPvrovSxpvjSXouzs/4pYx/ejiHS/O7DvUPxETiXvfk7
nxJXOqUFP/AdFsfcAxlmBT799UxGXqGxA6JZbR7WCMYvxLn1gGK9j8MiuR0IsAWAGOretaKX9VtG
Cfc7NZumPVM2sNyK1BbgDRYPUcFF2gSSL9Qd6JAfoRhxCTXApk5mkltESeMsUcAJD/zWgdzwIchi
FJ0SKgwfXeWesm9O8MlClj4afFrE6DJNQsp9dglDNNYTutYgVXH7psATsepxBuCw1IrfDQoV7xqM
IlZPtwnlwbIr2ckMCGebm6o/yxC6YUKKpiomq0/cwX5pczGYLIsHpkdHbteeKsvTN8oVztJh9ubI
E5eH3miFeDpTVusIpNfR/yElVINFZRQ5HXgCSjm7NCbyFEHl7d5JjW0Tf6kh8F5qv55JLofGxNhD
9NsAxxrPb6FHPrbWoh/ATOdn0+YCtTUBD8mPxj1iWSyp3XJrOGNAcW0ZMeQD8Jdfr1P3WzMe9iyO
sgRTf/uPDvLfkLL67x6gWNpROyXKmoLRpTbbbkiCdrf8rSyQWnKKBEB8essOKf3L0PPjtHVP1J+I
h01xvgZGoTE1WM4inwpV5TYO5ifT3vMfsfnS1TU+Q/vMC2lj+ye3DQuVybtiQmcgfNvWeZAH76hV
D0oTWaHN8sOafHMIsKU8zl0EdlAbc4pFyNsshJ1+IxCtl76OrfTJYlPjIhbGzMngM2Q5hC4pVWug
sxvC2QnT9+/hRY5SX3GKPFqSRdNf/aafaH7ZUVZGlgOIY12ALoozO2vxindeDWyJONRt6lHN0Od2
DgqPRa121B+nt7CTNrhvwRFIEZrW2HQkkHHs0ZOoL3XKcZi0+zQijgdTu6Aa2xMx0JN8C92OZKe6
a04DwvURdWkBiy46Ij2ocAXqjjsUiAZJgLK1H6Z7M24MD6V5lhqcY8IuJVRSqMrhuJRcewh2iWfk
0l9mT6ZFJPUT9iW7LtzWNpr0oMG+Lr65oDNPGsCS9XJQPU4cP1igUpfgGA7/0lJOSTaseejq//7V
hFLyeQrU8BZpgd6F69AfZBN6H6bsa3NvqHd8DcWKVnk0LS8pdUOzLoSfaJ7bAVxCSFW8p413vcyy
hVIor70D+tgyNJzd+IMNhws/srACaMrPW4MT60gIzQJoXGVP5qztkWOLvDR/7A4xmU9t4qHdREZp
tcfZnzvFNH3nY9zatiJ0U6AXDtxy2huXJfkcHjSau+WhqlE4stXVWAz4U/7H0VAJUbrTM+obz5Vi
/vWL4zajPdDx1bnmEzcvXzNYpKw77a05x7ZIHJl+P2etxoLSvOW+buHpicqm7/WpvO4AX3mZ8jrm
oHB9CoT0/fgoQp+O/ZKVrMKn/t+ToZEd8K7pGXhTYYO6XnuDcl1S4NeaQ9pv25vVli4CLgywLEEj
sWVmmy2dlMy5gXQh33hGOiIp6kJ76I6/gfuzjnXVCpZccSp8IUYC1+br2mjVxV00BOy4VYcA2CMc
PnLAna+AaKtMZbKPeqhkjRcq1GCBht07NQw8pMFzNKOtJL1pvaQo2Pg1xV7kbYmmaHc/uUrAO+Dr
PzHKNHNLjOIW9BoL5z68h8pNShgkrForQVYgx+xTHLTWlclBPSI+BCurIj/KzupCJ/267ctSXRAl
IgLGkX7iIiN/6XdyH1a2lM8fLnxyAKHQhUSb7KLh0o7cVWnlZI7Vc3bM3LthZIRT0r2YtAeLrxi9
dNddZ5amCGO7zM3wq3vRBo3g+DdPAfQ9hMHU8QmhRPFTVZdOczgQ6i5R4cPIDtODXosLz6wLmEr0
piJ/tTXeFuqB35WgHc3Ar8uKN/amLED/uGTgz7eHht7XoVfsxkeI6j0TFa+84IvbsJ5M3fCIGuhK
HhbDz0Ac4gigS2cIOnvOO7sbdUUAe5rd3qkaVMow9IiTGhHLhc0VSTF9hNSxVaS0u9ajivTXswcI
ICITJEyUeK+xEnvKpvNTSTYty5cwBY/lC4nV/ND471bnTaLcH8eDOfaDxtYmPw121RXd1Xsvmcos
zTdeBT+wvLZ0EamkqJ1C5M4yj/AxeuZMx0tIacgddYHuhL1Mx+G4Y+hWal73Zv/9Abz2hJWzfBBm
oyuOozeMj3F41X1PNR+vfTuRLR8SM7zGUAEbl77SiSpwtmFAD360NDgfKoAk/WQo9mA4JFZjwK4a
DoytaAfyECgcKks4gk94w3N/zbq6ZJmakcKsplg+pxqk++dNblQybv0bnjytRCnYxlC0Wn1TJDlt
2xv/kCWRG/0EiWVlSL83Kr5Z4LLSTUJmZb/2cJP0+8ifoUTv9aDbvjqPrf6u++a906I/joalbefT
0f1Sa3J09R2OflKr3IqFkvQsHhAwVpyKITDlMXxhIhIvm3u4kPxspfehKX9JgFeqNEmhbgX4bgZR
3RYL31+IDUt8MvsHEZCiLiwO4waARyAHwFbz8RtI8BmPyY6MxaY3IOyzD7jToGcN1kgghThqfQev
tOmm3RJ6LmDR1XMW+22u0sCnxoNMP6o+ve9SLrSKVitSoPsUDAsKIfFFrEGLysCixEX1pB6HLxzc
qNsuVlzvpsAy5TnhD+oHXVS7yOVesf0hJYTnVtIAZh550/fu7k3wBIIHgD+9x0COJhK5u5KFzk4/
6W1Nc4FCzwR5JDODXq7YyRuC8DBRE+BBlT/pX4faWUoXEY5kHI9zsPE8QQzDlXffCMtBJN5fP22I
n9N2nt/K5KVOlH7P9yMXaowFrMbdYazm7QgvvimrctFLCrDOeGaFPNZWSP3KOK+FBFnih9Ut5XO+
RNwXek+gK2Y1u2ijvfOf9FSIMDQySZIMuHJhZNq24Ob0KfNxyjobu0UV4AVM30NX3Ojl7nsB/Aht
EnIqz1UiQ6CEb5eHElzMv7i0w6Vy3RW9h75R2uMyqQqHH/tI+mjN1NQyFiO7p7FiDF3AZfckfOo7
Vgaf9z8/ThzlbIlJWHqXY9qdUKg2Kt1FEPgLxPpmzfoBXNCZp++UDwNdmw8m870xE0hRuv4HyXpQ
DRls3fK6q1Y3qQfKqBo4hFPIW9qRopwvleUDZaEyHMSikvE/MjArqrquyIPQPRbwP8XZFH5t0XNx
U514isgyBXGctS9D7iL7m3NCG/2/lfT3pCmw5JMQ5cy6yPs3yHjNcA9TKfDV7mdP+HnY24QV9MZF
wP523awlynfDoq0Eyl8YaMwggDeIg2rLbaY+DWh7n2Tur9DQIeXssT7jTQxkAlKa9xz0N0inZqqJ
Uz/1R+V8oNPfVWVO9/BArVno74y6x+8IJQMeACt2Gjfthxt6Lq0lmfylNl9fGOrwGvgO5vYd+rH7
3H1ga7L+L9AyLFV6ViJZv22+YBDJeFNVANRaM505YfjDoaXfNnZgET9ngvkaPd5Dg95qHqS8oISG
ozixNGaA1aUt6u62OxmjQN0spBvUedOL2JV+PRqR9hE/0N4aIJTP0r34G2dk9za6arrOy8KYTfhJ
w5stEroUAyb4+Zvb961+4ecDXlqMJ70MOPIUnV+Qi7Atsz5nSd//K1Cny2vzUsEdlbrsEASGSHPN
QYw6N7nBy2GAGkPkvZoJUz3XSGrrClIF7oFyiQBi+hTohEYuG0r/3P0/7I2icceWZ57LL5bhVPxY
/KEB+8lAYVwhuOV4p/DzO4phQq9w+o1UtmSp7QkUkZVRR1EW64LGjn21lxlRCg7ghr2r8Aa3gl4W
i9KWfjL/faese3ku2eeW/6d+AgJ43bUAFLDIJ0rDRNiuErOotCqUByoftUgMDH9qmKyEHk6OT4Vg
s2d6Mbz7k2fBC7eS3l43Q5968gCpNT30W6kscyLhLMYm9k5+iZK6+iY5xPkmuMkJoBmiyke/tg+w
VuOPX/ujAYDZg/qTzpZQ7RIbqSWoT2V4x3r2sPpEFgjQq/rrr5k2QF/QFy87K7vTWf9WPoaEK3YH
uzYuKmd3eyPH+SfEZrW4L+jomknndG67aPsPrT3wAqjYIxNnXhyu7JRE4cY2SbFKAAiaHoEp0H1W
EdlF6lb2DQLqdaslj1aDwRom5S/QPoc4iHr5tzf4zR/T913CS/X6bsbEfSXliaQ6bNw5dF5vauTC
KmqhTFNaziEBiX+xfvPKwKU4lhmXDr09u5yBWoYrKjDZ26DgIVG273sEO9C30Egv/upHooqE739k
T/+1XH7s1AlTrky9WlktO6KV3Ei6qfHLfSGhkXVH7s8VwRaJxJDZQtuC68E0CyRxF9ixsevTtHTN
re0sK8h20iQwnrSmavzeMd6FlniOneMq/6yP2/u3Z3gDIJotqZ91AsC4dg1AttRN+C0mu172B+q2
x4LSnMyUJ1nZRNNMLHVREfRNF5ZYdKGMRY9eG5GYYof8x2qon1I4VJZuFOnaeudqZED1ocV5d9wD
H4seKdK7Zymf1zT7+1E2Tpp/a51z5+o5N1fi+uPMuliPzZFLdF2Tnw7+SGD1Dw5NM3COynydCkJx
jLs7d5vmuENjrNnI7ybat5hPb2luld3rpP2x5sLgT/6uf0de/UbMtuU5duTJ1oDo4fKzhU1EApLq
rnI69aIlyyH5b9qNnc1hE20FCX8uhAFTvXrP/VrVlF47SHu+lL2O2iT1dcX/8aWbmRoXUGrM2Swe
OsccwAnlaSAUUwcp2IjNEwXFv0OCA8WxDYmw+mbc8KaAME9ZK2bKaOTaW7Zf8Qpo3ScaiZziBcYW
i+Bhc6YXbW0iQAW15J8VRMQKpKom4G+/bCU+qyJWW/5jKsy7ZZ/cuR3frviUJU8C3N9ra1riVCbZ
1cEXnYTV7PwoGW08FRkJlewafuFtz+hbvGhiItijbd0op0YVxFs454/WM6Amevc2/dZATXKiP+jk
wFwxf3yAEu+Er+1sEvmCg1C2f8tBllLm1sR+HILVY86nKGth88kP5Jb4ryYuX86zKcetfrPBnYQz
+ksbNUbv7uE+BTo0VGPgcw0LEsZlwIe29MYJMatdXI+B/2xZCxdHFeBiHn9tAZTzbpox6Mq9PAHF
FA6btCYIewJx5Gh0buewMSjFiIKVKqSGg7Iql9FT0lPulaMm8DrZRLXkg2w2epiXTDbgZpkKRqq9
0n8w+AjDp8hIUsV+5N8u8fZGk9tN4KGdG6DObvaMXVnYn+gjo9s8/AiULTVblPJ5o4YKoE8UuHYn
EI/uVvQW0B/x42kGugSEjqolMMFXtUJaCb+FoohhkRXFqF5JMpNbAg7MXA8pbt0HUf7olDbMPT2V
4/cTbjzbHcXIXwEg17DWXfmhkt+Oil7Jxv4mFHh1QlKMprC7UQEkXKFCOHeLzsc+uI9z6PUYpK/7
xWweqTJwBx18iuZlUezRaVkHQ7/fDb+oS8hfW7TnBQhbJ2m3wADR8wzmYCCMkZmrAAf1QCnzvyMk
IWkya3+AOW7p3joTqWf7LFiaoWvV/zJKY2zfkjFbGpMJ7ItQn+DuitQ/SLKyZjNkoRZPGI/HI1u4
9/vOEzy4f4EZm1+bkokJL0VL0qUB0GazSIfiAMqwrlpTE11R+IFMJHBdCJqsVqjRfaqimmT+BXlx
b2fiCK8S02FnaHUwg8LUKKiptkQrZQQDQJlspN4DI61zF7WifczPO0x4aIt94h5TwdGW6D4YvX3D
CvM3xOHs/8UDR+e8qYIvJXhlSRxh/CnB+xcORitQscbkk34pIOYjhbLFNTgXDPhfL4oD4Pz5zBaf
aCCyfhojqlHq7zEZeHDTpFccH5CHZEkqoklErcqd+C9NcAutIg/navOvdGwRVvu4Gduhdt/zkVmB
c9CBLBpUyk/A9EKRLGbq0ODshrdrs/eoMm1w8BKHg/2cAlxDT3SpikE7UpVMz5XKXiCYzIQZHc1e
meHTL4ftHL4mOD9KmF9Q70reu5cQtfN9Q1HDtl0LNw4lW7h5YPrghEXrJKVK5ndcVmKSiNv08VXp
OnwkoZKeJCcIWpE0mvfGjdO/QzO8Wkhu8zqaOnU6hk65ESDPH2KMAbmSAEQiXBgg+Phutpru/EDW
UXxQWmdkjkXWwqHINWLibjU16KhM2OhLnS8FYlVxRXoCwW5yxlDPTx09zDzPeqWZq4FFO0N+nUEV
M7zyaOquAtr/Zjc4o/ZBktYxUGUxaE+MZGMqEDdP9YwQezxlrmLMR4xDJWIKhryiCjhF+7WcTFmp
7HqKv2u8FteY2esGz3PtTjZesBMfCf1j1EjVXeEPXT2CEKv4CttlOUd04v0K4wjtXCAdhOV+PS3r
eKadahxWxG+XO6uEmFczwu/PVIKW2clb+z4I9lfTHOYTXFs4iruoaXoJgNOmrFf76kPi4VKUAiDl
7G9YRpV8nQvDuxCQc4ImPEQe/fUs8vU7GI6802CX9yhl3Vh4Zw2MPD9/SwwolMParx5rbYkpInS6
vuEO0iJwQJeHOhm7inbFVUiX3wlEJQtbWt/nArFKR9ICyAt4P1maArKgmKLS/n3EZESZZXOuNfw0
mnF9Q1g+yTL8XNAC5VnKgu/6U2wPlv6PFbk4wmOx83H9jdejA9mQ0/wu7Oxrop81OCcO0mXMb2AC
bINpBMBA3TtLYCQFwhqVrOtqu1sYeh7vXdWa+xiNhPKlnRcFfQ7APJM9NBcdAh3X+3mYOR8dOnjK
cKF9egatoHbJbhaXBoIS3r8MlS5FYgK5Aotk36zi9wgQ6VKnvKLlwfUZZTmiclAIPi0B0Welo0W4
MuBoawI9ElHX/QRhJ1kjg8t9R8qlal6jjQjIKusycWVrGd/j+H/JR6TVlS5O/kLvRCuljRRBx+Fq
rjgZ40spyLp0KhWF0e4FiTitp3yL88m9LuiH5n9vhhZsdD0JvW/Bpkg12NdWQFTFImBWMmaIoCzK
kmlb4xFSO9hAgr+GBnKRunvaNwkagXJnmbm8knP7LFsmnpo/TumMM7Ubj9Qy46TmN2dWDplZJrm/
ueuTwrlq0RajGI7tmvcqY+MEAJE0HkCMQznkDTkBXpOqMW0y9WwFL+JUDUDHmcGGEehct1vPPfOj
8Iy1ZIViQ8xxlVPTugwzi7c8nNHgh7pFeMO17ad5zGDcz11YtSjfbFO35ZdbOLjdrdj2ODMZxtci
CesTWz1qH0WMjeMPGSSA/tOsatGUMaBkmDrUxYFGmYU6MqmWp5lP+XXgItjRCST3M67ot+nMyT6T
mn8Pyw5fm2ldbwaxfNUf5aGA6wzDeyaZc267l2UK5sfd5W5MISJ8cRFahOppR6YpmxfQMK+ghknk
RENznyKKMRgrWZo9Qt7praIFDYwpQfzD9SF+Nx6mA+AnwLFZaqSIDXNY5YPnjn3xhn0CN1ECRzkK
9bXu6N4Jpl4rqfj5dpsX6KbDGyrPMm74enuu0UTezj5wWuqO8ITOJSE+OmF1woYNwcUD+Fs2i7Ro
YE6get9vX0tV0jANbiVG7gEqgNGf8Ax/PFPawidH9y5dhTZmdXsw3CBXOv64uMjJjPZmdBh98XqF
7iR1qooe7kl8SWyUsxfZiKMM7YhBShHyOw2wNuezwhGTtBEJO4EHU5QaVF9MeiQUnOuW+7XgY4Y4
ZIp17sHRGh4u77zJM1HhOVuqlVtVSUGPYgM7jaYE1cj6qGx524xHVmy+MpPLvGrXUmxpntIs6D3Z
TUOLH4LzImMxLVb1GlV2TW+J/mmLcZLgKP/P+g+8EKetBHk8e5y6v63V8zqTEzxdnWXMjZfowXly
7yRTyGtK56I+4UAKzX7VHhl4tBNGPuUJi1EeUpvM5oHIlPp59en0UNYlsb0u4iwzkr59DRaqAGei
o3JPwzsgBR/bDSLKahBtop76hTvAtlYFfxkYVU9LNlI5EksYM9IOCGdJyUTnwUKhj7UlLLh9ydMO
Va7RW8sRR7MTXrBzXcElCh24DLlQ5JCnyjpMT6Xm3Ypq408suHP0JC6BD8Cl4uP1QUv4dP0GNzdX
JVc+IToevEogmCA7cXw0//Ab47GmkEkzbk3uzbqlNO/4M5ssQIUUK258FHjoZaFlK/2xoapCzMn5
M2Nrs19KGtL2e+CzroxMfyNtD+Oe9+RLmuqgSKnuvdyw9epqsdiQU7Ztm4+qzL7jMJS5awC+isNq
j5gZ+O0RxusgpgVT/9TagbLJrPwSZictxGvf2jEjuie1NUo1cxc/xVg5Zh9s/Lv/D0qiAL/4SBf9
Kv7XezccH13LqTSp0xqjgtZUnZ7B4EQ78/2ZaeDE4YJEjLdqW1JcfvkltkYjhqF619MbtNeuDlvc
NFdjVbs8DXkQVR7CXwcFrwBBK2ozoYOGQR8sMacHQ3B+dqpncMWme4FqXTYMeu2BP1Me8Ot97R24
SHZ4Of3ZCuoz1sPwG0vKqcFnqPMKC+/+1Gb5fHYueQnjTHmSCyAWkKctqmyLQl9z1Hkz1gKDqYti
XIzRx1HPtgv7SAFfVEWcqc3kOtvLgi1QoGNOIpMLlOY0h/qdUo/Yshwx8/b83LLfjcLxPadOQ7X/
mpPV7/cTznECdyxyBo3aB2pMQp0AASHZYUgGMb8bk8UWSZ3NXKvofELlrxfvpWRNygNWRFjPgrjN
Y2SfuDp9975XUqueB6nTqU547tJtM25s6mjoMyDX5yPYY8vy+zwrPqf/EEh68+JB82+c/lo9MvzY
m4uwU+pEWga9gTfxSau6co9y5gwoS8YSXwQsCIKlOQotAZHTf+A6LKnQ9jlgQA1Fe+M4RjpTfBsc
jykKdrfdJ6bVaJgM1UNhfTCP3Z+DEbSTcmwZiwv02IsmHev/FBGLHhyN0PZtlzF0KH5NaDiQQfNC
lckXvzVAliC3PLO30G2SYf7x0y2+8w/7mMh5uFaWC0DtXkPsiaEzfjlH4UBXulWiU+f/5jEOuY7l
6IiW6deL80IGNfduSSo10FoGqhSqglfGHjq63my+HCotPmXuwFA04zzfN0X3QDAGAEwcIuehDPCl
ET7miaHQuDBVJekcIHMdYXWV8sOfGAGDMo75Bkm5EY1fs73h3FA9Sn/gUQz1oFOQLbPfRn+eaPUW
MDJ3P5k2tKqa/OjRSK0qG00tZaOYcwhmX1LfbXBEeIw6zPNn0VAxuyzQXMMiL3PuLVaprou1MK4h
idEJSA8PVthuAQv4Sgwo4gi+1L1YI2fwd6AqtVCBfls4/lI2UWNZj9Mbx4YkUvF1GZA3t4iqHeR6
+ttb5f0aCI0oUK3tVNTaHxeQTf7MqKhLHSgvGJ3leymOKleij3IqIIyjdDaQahjYVigbX0rTFQVI
en9Yc9p59mHL4Z5TOEHoXXPz7y/JkF9Ry9KHjhc4ocpSM+nU7hka8r7JBVd7HtOtkf9ysLXYxJ+Z
sB17U+1B1HwQjwmNX9WIwl9Bf+nH3gFoeth52zbqJn/mTIZqOH9WofPX5M7lfw2Hy/yPZAOtIwjB
HhQPS3DALVbyaydHyM+iqXB3dwnxW/TTM8FYs7wm45H27EyriOvjS2oNF9/MXZxPfsRXc0qCCYy/
pxumZ7lpiJeQbWt0lse/eLPe+rRbuSWr10REMeH5Rv/xBR21c+p+pl4a0sCKSLxRpMFpukR6tv//
B/XMg8ZlmBct14GJ46BJfvHuvA42y6GG7uAhOR3gILF4OvTzZQIeTqTTG8VK/q/V8yWGGt8xTjXG
nEPPan0RmRneAmfbuu78HyxHZ34+EOUrFrYveYd2s3EQ9PcrWGxag9j0btX7IesjtoM6YHkmtVXz
lKx6uMrXKUb0qFt9r9cXdFD9V7IA3djvrGg3I1skEKL1eN+zEdyHDEXdLNGTOMBf4Po7uXexqKUr
t5IoUnHXjYkpyaDBqJroHMiyAUh7Wnct48rnOF3JnuEwP7QNdv+QeD/xJMp5MthsRvnASEqKqYJG
u6UhHabf4pJuskwOLEFwo9MlHls1jf2HBW01JnOivit8WCHb411m/u1louL0amq4GWLedMttcsoK
LXZEYj0hRXpV8/3cpccJPkVGJqrRMeETGmBzsnf69eG/U4aO/SqNVZ0Jt6TgTGTW58+HdA//8Ktf
AaCvdmDYWShcKC8zWc3CsN7mImJpiRi9cJfy3W7G/CFJrzaXLG9RKejdZwe0jUPgNHF6Z62JZwcW
tmT+i6egFqIC9Uf6vowR4RYz+GeNmc4Nu1/psK8glFFhOfSsEZCVCyOtYTT40GPEsCbOTHH8DEmk
n2Ad5nh94yl7Yt0QytIW2LYFfDdFW/q/HSFDrg0+KDLd0aHqykSCM7cDnzqJN72Y5CHxXF1Szdfq
yb2jZCEntufIuPH3qsMFwcyfG6Jjbdpnqv/YJeEdPoWFjnSBhre2ApiS9nM+Pcgqs0bDCssMMRz5
yh8fe1kG7L3a98rHBSDm9fV/Kx8ZDXSW3TShShsaNs8STIu4Jg3tGqX2ffqiarCh0KlAbmDhLirr
QV6m/t1allLe87IXZyd1jG7mCK3g0/p5ERsxyUP+a/vtixMiFzmfDphtb0tyI2mw4axTTiRKm3HD
5bdDjp4xSRUUqN0urHxEQSJL8ED+4SlpovJMo31+YkUjqgXfIzLXIlb1dWDSCfBPGgKaHjeOLylV
onT71s2F3tZMt8M5ZBd124yZ7GKElKNpcpPJ/X41+O3AfgV9Ev/fp+c7ZfaAngy497b8QQoJZWeV
V57QhFSuehz/e4mQKJ8lc1ixIZKXARkXHQn9zwNCyMpdYarc2/NsBHQyPS+shG8RO/CLZt4CIixg
cGSrD5LNCEomluwv9ImSqt5NmiuBG12/PGEJRjyug4LeuNEIbIsIQiSP1uTyZF65sxQK3rZ4OEMn
nEBT+caZbOK53oZj0YM+Y27lM3ah1ASX91iLKITT1nGlIYElYR6sklExv4EsByVZIoc5n2baNKVz
cXGLUB0nvjMQqA2BfE18AmtnFtMx1tL9Q/w6m0z2oe72jinKrOXwC52I+m4FmEvQpOMCHV5pPih1
KigMsJijguQT0lRQLxpHR9PrjF4ZTt9p3VsXfi8QseBkLnZGCsqGOSQico2pkfAPbZ9ynaO1IAZw
dh+zFv1LHElLshK8fuXTpNySBD5P6osQNdDFpqkXsOHKZSrobPdxZn9HzMZIyQhM5YkWXpcR/Pi8
o3nVYaBMHGaV/wNBUqvOBVxTH4herx8ddD8MjwBEKBfhFq9GzxybY7CWUMZIKPldkj/57Bywgasg
BEL25iWdlod29qTa4aB/FZ0GU/4DUse7EjixE8+a/rDbchFw4I6Ty+hSi4d3+tGqt3D6sDlgTeeD
WhGJNifJl8OtfgW3eOdn9+1+eov+dZgkI1hhdB6qav1+dbJQgSd9f4snauashZ1Xi2+IgA9ci/XG
61/oyZyMeCSz0YMi3RQLESXi9UNRmSk0CYDnnAWggGdvXeMdA+cVAWA0sfPA2qCIJS3Xi042xlr7
rGhcQkbqUNPUx2WYxyD5esSmB0d+S1GoPhCbcKb32Ri+ITVtiDYsGDlnbW3pWAjnhhO8HYE/Ngfb
sCsTIM4b8R3ihAh0qJqFa9pOgFBjadp+mygq1VjQpjvui89AljttjkBAUUV13gz3A06mxKhEzEn4
uyjziDWboGvTR6mHhAd2LC/cw9a0jWLqUQ3k7YUwOhp6E2rWN0vJTyP9w57xwmoEbvyKmfhA/8oe
DVi1eA8PrHSyftLlzkvtQEpXXblfPITbniLsNwcNIDn53xHNLSTo/LDCUZF0+S2uG/Rw0ZdIi+YO
djeHqRNOxXEz8gWtDgPasYDkrC49hpWQRv7gIlshIYd9Ll7Lq0ax6dvZLHnwkGcz5EZ3jKBP1eB8
Bzc5lREGRP1+FBocuS+HW1uz1KIT0rWEm0X3qEFcn1tHIjFEbhmfFpL+7XZZF1Es5d9o4xTpukKR
fA/ntt5hX4GG4+AQcivR8ctE+14Q1Kbub7gr++khTZ3yF88WUt+RaEUCaR8vZ7e8pq7AUopFysB2
yAd6m3yrbcsG/SE3NH0j9YIuTHdWj061cbra9ZZ3DIvkO4kIMN11fNXd+7aaFen1BlotfJXKAnfx
T3GquUGkxF8u1+j5lFVi2/YDwzNbqQMAC1Te8Qfeeq5lzyuRnkqPO8773q5p3u/H7Tyb3dF7Az/f
SUop3E5kjaSe2V+pyW3PzuxyDVCWkJnrYMRF3ZCwMz4L0NTNoSpyuSHjD/V5cYhNnDlpThry01K8
A6TmeIIB6CiirwhwyyYh+B6r0vZML5u0TjbKgogTw6spixfqNrJRjt0njSXrxfXJqk7c9soywx5c
kNWV/CfUchDzkkpCeLzcvuyr9XAMokr5B6cR0nL88egEPoimiLGUUubPo/1YzblhH++msStVUqKy
RRQn+h9qVYWlTAO2nXNN8yuw2+5olk53cWKjtLHw2cqc4uZ9GyL6/PDDJ0fSWN/qfFJqfBgv+8dh
A4qr76myML3ZvDshSjXrl41TRXbA59eoIoUsY/6hhf0mx8Nbe/7MyBTR1oy8KGPObmszZB1K3vA3
LX0/JoLTAmiKKuRtH8Md3IRA1zrE9orDvGM90BydkATKa8VhfortT/Z/ltPIOgBrAXINEpUn26Me
lCN+Nw0sN/ZXLK/9lrpp9cLKDA8IHxUdEyHW7B7QYRUPGJjbeEqCxFA+Z2n2IcB/44xwDsttOBon
xtHZkxVfXCdBhTPUl0mP9RPWGrx8VVOFI4lbJnU0CIXfHHHKGObxL1iYrW0gNUT0sDJBlbtHIu14
Ih4LfWJt9VF8L135we+kLWkhL+Y5mXGar/IUbDiEI3RxvJyg3Hqd7F3qHFjoDXHPMef70jzaRY48
TKBF9LdR6vqKStITAv3nPG8q4Fjr6qb5AajoH4NLK9aDwkCFttMUsofi7Zt5jCovbkmm7AAsO9Oj
p1jgwe9yK1kCZB3Tr7t49vMcMP0poSGCXnihPLCpfskPoe9WCI5rIWR07iaLPKimcBskDML88ucn
0H+qHFttVDZU/YGK7V1Fwx8WwQHpdPPZLnbbEuwn3fK751Xr/uSlLuQ/NEE52rqCf7xKwBx7AEjY
CX1PoYAoZeyg65O4XZ+WcOUl9anXUva9gNbLOxhYDcAPaKiIMczXq3nEQ8xyYpnyNpriwBTUvn6x
6+B8+3v/jlqIMb7dY+0L2w+H8119It3C/2nJwSex/n6Rswh7QvStzKLdqzcyX+kpwXxbTqv8Od4v
GEkiml4q9iAoReODMh8atn329d9gePBqv/5FEH3igIaYsNHZhOdQ+m9akhCuvAiKr59uj0Vhg431
cn468GVyua7KccIG+vglVwhBK56sAhk/WTzBurSyCMuuOnodle9iYX6DFo83VhC8lO5VJwDuTh5K
EZVXA/two6dsIutYnwvLt9RaaPA/I1dTA4G40xmkO6N3Nh9nDJzhf1J6iH1MizdNwtUmkgHVmxB5
jryIOoV/qoPi6vSn+pC7fDmhkisP2ORH2InXhcZDBIekQSRdz8Qn0GRvtEfD9qbWHGNmXcm6d7F2
ckkDfYNdzNm5UoftYK/MhNqMJkEKLHsXxt36941/+sdnZVr1oJRPUuEaYp5QkdTFOvc34GwRvVlQ
8WVY9laZcAxvlqv/PtCVbh9qeB/WiaiuVfKl0Gh2KiDUVrTUFDEEWHETn1hfqFJCKxiOUyLHoiWE
GJWtTYKcm0Qjce7nd5AzfNmJR7n5u7ntp2zbh3lrBDDBMbS3r5JLt8PhHKWsSnGEegRO5t2JiYGC
Hx3XvNSDdj3YkVNnxug/Njrb8hJ2WEpnkZR+tF41lkeR/CuBqHdHw2C4ePtvlOm4Y5iIqxX/MOKm
Ar4P23Y+F7+Mqd27tVOtPZanbHjSwSDPB88nTLjyuHmADhCRHi2kU+a3+YIhX2PMkE5cANjKciW7
a3l60Jxyf88TZb15ipKLlyc7xAiDvXNgb7DgVH/CkWzwysdQNESYDrbacZV+XhudJ+BDPHZlMN1x
8pa44nAR/iCYNo7VSQkwt7OKYebhFtwvMtm5D/8Gm2DEN4GRnoHQTPUSgIRafxA9x1Y2iq/dTb6w
onlbs61jfd4g8qvoG4xaJWVtKPnvw87tD0DHrRNjOagAr8MXkzI6eBYAdcF3gMTO7V54jigScWIe
6mXxap/ZvRcXZj3oUN1uvrD2LzfEykrhoG6KdD4/YcJumrGVSNaycwCC93w/41mITsqvUK1EnUu3
JjwkS/mYFeZ3FQYsoX+Lcilo1VhUq2XZ9iNJ9bpulqxACeph+dQuazMUblnGLcT5YMriIzrJTM4L
TXsCJOjcXWwqMefdeeWXGPo9fVJyBZKkbTULxEtbeBAggm+eoW5QL/KKbPgCBnWOqLLtHm0Fx6IW
KyLPhlrLFH0dXFIIts4aXSBk6bRz3fbybXVz28lMpKIBVVozDpnzx39rcYccgwpLYVJC5vvDiOWc
6lF68yrp54RMocRJD62xBAMIAUu8HAE9OZgbRrq/fAl1cBgZgI0OeRtAowbfCxPl/W/mwzJQdIHC
VCuRx7Iot07SJFyrxil20hMr8QRmPKlt3Ks28a6ooFLnEEMEgWGM6hk+sgpiD3e/p1rJovkeytWC
CzPLDAUnQnI8SblQyXam70AB9PWO97f9s1gkm9+JT43ICEaZKQGBdzwngsz/3BKpzSeENOYjH/Dp
EVkH9oVWfsC0awcvbyjoF6dfbApX+3SmthN/mcRkf7GFn8+/O5nQEm1jrlUCcgSNY3e19iPC1Qlj
clmsntFFoKwOd50fBtixFiAUKB9hNo6fw6b2GTcXmFtph+DqX4OOHKwkcdZTF5vGi+UiQfELaMOQ
Rkd8OFHmZfYmZgD7feeyrLbSYwGgw82eW45IMmJu54tfqRONU99OPsoTmTYToJIfB8oDwDHhR0Hm
Ak3hmFF5dXqtfCqodqUdLp3aLStl6/Jn/NYNiuGul8b16uQSnsUGVjIA9FQA8JSGuH8VK+DZEMJJ
DxIGUI1E1Fwdtzrzh9qbp0VTtzm8bTbLfH//JCjOcKjpdiTpnVJ1DtGHTjHznuOJh0xvwoezuUOc
sQS+0V5YA5VNgxoDPX7U+foC550O5+NwnRf9hkAta6h3I3wtYStWNWRmSje7I+cV02YjgVh2eMWX
5+ON/DLaLAGINWKFumuBU1EdwNx4cQYZ0PTxSeCPF7GPdN/x1BKZXFIcnmiwbP2PlumQ37R9IMyo
d7ibb05pLJlDShMrCKVSkFioEBSsO3R+OZvJTrysdHImAjlDWqfkj6thmrWuEjF0lrEpdJvt+OKX
xtYfHOCnMO1HQDE9E6wVAX/So+j6BaoM540EzPP02rjB68C9B112By/5f6eKYVdaVVuJhhIx6PDc
QRzTHWZZGsv7HJDw/Ar3Ui/7pnqPMDeZB9WjZniyb69QTvbClFwrFZ227ttrJuv6Vt//4Hvv3UJj
ERhtGWkjKtouyur+IquDAnKjWx1j7849IVOacwUxnTrsXWTZUSfn0tmt0yX/CIfQzQt4t/XAoHKU
GHlEUJCB5DtVTYlBQApcQkxzD3y6GCXXYE3n5ZgFSBG6kpHtOf0zfxGHFKBWyEG4/x6xNs0T81I3
3QB1o2eQXOk+tHwwzverozQcjV5Z1f6lyXyIx76ERYffZ/zPI/WdN7WH965r12R+3wesx70EJEvy
CPDu8Y0/geE6RNrvaS98JXpeq+WPZPvyZ6IrnjfE8rKTBFDGVbf1NfhcM+KJhH4WJyGs7OF+0eNt
xM/Y+lOM4nsmhIH/zuScFYgVYXeXJv0vDofkZVhIo6Act9nARxsWvukizj2opzQKDH1mBd+aoWNb
AnqOpq6RIo8yAjeVO/z9QkelGcu6qUDjjwEzy4vaGUYGSmWSeGnVq0qwKKzZbPaxjESnY+Zuqo8u
yiLEZLnYc+sge0WhZYwNKwwVfGBV/La0p14ETNgCTfFWqfOI70Wfg+KdTSPbVfZyts7iBy6buwoh
D9H26SvZO5ce5K1zhcLxlj0rUtS0NtwE4BXY0mF/l4qT4/YMR8ZDiVGRTQE1+tl2nekQJtIoIn3o
3DEGhbTT/yRkfhYOyMCWoWhpDheS215uIP0p5d7B3Xk+o+CNQCV9TK1ZQRUqqcR6ke2R2rIq2SGu
Hwa/M3IbFE80mWanQAhkTBKJQ47Cqfqw7Zx4JyKR9MB01eIVEQ+1X667A+R+tlMvW+O+pJh5yj9N
wD9cVBDwZcTHy4qAa7MArsAqUYGOtb1/Sz5OPwCc/8UJEaWFqPm7E+oroKFK4djLPbfr3ieNMzBw
XJcCaK0q+79m8efh6CK2Z5Hl266I9ECCoIxDYP2jToJYXburqWNVH6Dgtmb78Z22JB+I8iXbAjfM
a6TTfTVxs9SrHajl/A6fXcP8Dd+LCdg47Kd6dgEW+F42Z9ebMR28xveuq/h3jQhvpv5mGURabIib
IBvyCexd4thNNEsLlDDnBhHEtjpUkyAVPURnvfoGNMswTc3jd2ACUkpYsWy+pH7josoRLnFDuNO5
LZIVa4qvAnAf6rAPy9Y2/5D4KTceWBMM89GQguJFiL5KXqfohZOXTMLpubD/Zcf/vazmj37uitkJ
0X+l8qIgPyLc2PTxhCQKaBZjn+tOVBOs6D6zlISpvuDfehNAelczIoM4UyPY8apfKmhxzL/wkbAk
rP0eCKw0EM3rhAOxh7h35mwGcdnW6G/ESRGoESztgwdm85AmXg+dzFPivLWJFyvOWnFlZuGrLzVz
nFK7QIAZeCA/KLPuaSJ7ZpG3WbEe+ZVWk+zxFqXI0QIlT7FvDAp9Iax2BsjNGHofR7lQrabUD5hH
BQgS1e2u6Qcyxmc1Q2gbvkdalOZOBvqT8xfzwVjS1rSS2nfo65hgR1YKxUu5f5kW0f9Gpi6PGSDA
adZA63RgI9IY+q5HpGn9zTo4UTRJyJePljJZbpZDzW9SGamZAYqFsW+NyzvWkGouko6tuP0m5P9p
LkJ4BCYyH6b0uyMllkzL/o19EfdJBTbabZKDz5b2K2EV9NgYjAgC9ji9C4ar23bizdnZ+LTrYc62
7iQM3TcxXLx+BmS+Or0M5SxSEuTPM7NQLJoSUSyWgCaRVIyTa/uZh1h0KPyqxkjACGc0V500knIt
Hcll9YLTTc3j1emloJmFJ68UHIwuXuT47d7mCkEkBt1TTzSCxYbQ3Ltov/m/C4qdA1J2Iy5/eaDz
UXkz+1ctuRxRXISttrIQdyhfvs+exsLHYFCQsxwPld3T0vaP7PiCe0/wkkNRlU5yafKulmNQx+1S
m8Uf0ZAD5wCuc4ycWk+HCZt1LsyB/LEvXO1TokJxvi3SG3n/IQHtPigh9td/cjYWiYhkU1JQh0ha
mnIIQvP+ZZM57Ca0BwjkG4sPqWU5qpfy796G3gr8+C+SkFq81iciKu4dbfYKOwYn+Z5AKKE2QtkD
4Ggh042xlH8thDoZP8H50fr2Sp5o1v7vJdmQWqWTNavamFp8WqzIUUdjWSjxgpnPGnW5WkokWVTZ
x4HU/TSTT2GVM1wx25YS/5FuDx9d46+XyWY4y3WjxFlQ8IogJg+KUa9Ba0opLQmBFJkB8Io/9+i/
NTtqBl9CM87aaFtb7ZJUCzl8i3yr4zJNLK7Xolg8eLaBSIUFteoq5alC73psROlJWllQyM53yIwE
VrcHNbOWGS8OWaYak4JTZn4YhwYXedgAHmKNJNlOjJQXHEDmYSdnUAmRhhEUxEYUPCXGsX+uQEY2
LrPbnT4liBq2ysyzRn7JGFpm7bsbUe06KgshD9tDeLhVYPTnMpCPknTogktbbH0DTuCnlts8b+Wv
7Af8PopcyE4LEgH/AwpuzhFo20RY+CWkSJvM3R7qZpeRpiX7Q7bviX8AjhkLRzQzMI07gCc1VsF6
s4tUkH8AjcVF6ZZrEUq0QYdj8PBoHu/6/ZhNlWKzOrjtMVopdQl7ZJcBmU3xfhUAfI9GkhwUHZdw
yq7lVfhNUngNJMF8aT9tl3yP419wDHlSXHbju4Oi+4auk6+p2GboQeReOaTZw9KoAWBZPuofT6av
eSzpJ2u0UOPhKsL6nQPrpyODmVSDiIE5nBUYxl1qnfJIMUf7LvAZ4t3/SU6T5YGto9/U7tBcwbr2
VrLr3GvjfXKQorEeKYZIFTbB8rkaP/abei1cco8sFwjhh695oym5qB2CTw56ZtU7NwFkSsKQwRQw
F5N2J0XN8oQJubvyxPtdxiaY+EjyyUoM35nAT4jjY81VYpcW6KAzpNy4dxxxSxY2P0e2FmvPd5+Q
NX8DbcD2zyU5AdZvDCYtqoosBpy2vZ4BTwsylI/CXpwci/Tg0EBNUR6M/LCoFrlvkV7YWIgeO+x4
KvUCbq53CwwRBvaUYlukJ19SwoaXI2hUdzHCU9/E7ue/BZLiphcT5IWAub5CqbaNP1koFPO8s73b
vLkciSq4phCxLH60Ze1kTB+hNxWlkFy9lCDoCvDbRtodXDlsmmG5GS3PJGByG1R9XJM2J5swTva8
bzlqX3hUn8uhz3Dj2Ka/bto3XJ4EnBnO+GFGiGpBjgsl2YqyDkSfTgqrDFqNRrdDwg9th3sDx4/u
i2g3rRVjn/x8piv7KC5S5qekcTwuV6P6xeis3Z1TbKF/ki393K36CIaZk+LtDutq+CfRucmnJfK5
1FhWv3b06ppQV4E5rHlzXo10VRgpRdEeKV/bTeHEMbUK3aRsJ2B4WkIlOh5j+lgoGa3+CrdDJA0I
uE8t+IUQZghGX5sBz6LdvxxSbgz3Pldivc3ba2aGGYSju1Zpzq22jyVsF3TEWTMtGGeXTqsXQCyz
bbkqbKd2ENDi/fiLL0ZK4TlbdMqKcbRnsvOVfz8tSDpUoQILaZ5ZyAu+EWIGIKJp6lr4oFVjUr+m
ldJclALiHQn7BvHCRaQTo9jnF86JqvtFs3xmXWwSs61xnWcO4Q1vcI1kI+yB2oE6qQVklt8u9k/t
raG7qRGLM5Mwl6DK+HBOAItDN0kcTlbk7xfWeO7JUO8ZFmoY4blT/jwWPmscfA48iTNqH2Wl8qO9
4X1oNyeN22GOmcqFrF0gU+utG38WwN4vhaZn7Fl09OHQy5yRxmxTOUNXwYT769bGpavNLiAZXHy6
CzONK0vFG8nn8NTJf8BDnNQ2fW13IXLDSKKkxKyT7CqrXhpd1rHLuwj4b80I4eKH//k0ZU2EbF+Q
joxTu6XSVwkH1pNuW5G++Q4Gf8zc+N8qFOIIHZiaXNuS5C9SSh+iKHP+JJMC0VH91Bf25Sn/ovjE
or8a0vqeOmQEaYB1wuz7P3UZtR90hekZNQmHFS9po+O2xFLunuT3FLxiv7vSQ94F6lO2F8petv7o
x9kBTmgE4bpCZ6WxXcPSHwoYE7daB5KzeTIq2yZSBCE6izB3m3cmo32R2TLXED6THp8e6aOyVeNA
dzpc/jhn8Z74nPDmiVkbZ/QV9eRUpBIDk8OWwr2dWxmP5EWRm6geEaboRxXFS9myA/L3Ud4Qc74/
Vxxq3lWIFLeWNZZvp5Abdp+YvSaD3EzLPgvl+qXeFmqXjlXJBpYIF6LYu2qkCFgTSQfwJjFwITXk
2PC6wbtRX9dQFNNjW1fcv8abMACWZ1hKqexEtKFoLqG8/NwJ/LS0i7Y5FQrs1sbgc43qniCW5ICr
u74PnptFQVlkh+P6Lp1kK+tff5qoqD5VACQ702rQKx6VqRh3Glk5cn1eQF+6ZHIuoUXjHVVQCE02
eN+jeIeQFWqRkcJmHqdF0GPKnXN5fxB2MMrgR1ikM2gNKoBhWA/aI9aFNUHmoLehEPV1rtXaczyh
GIa8y/2NQNlmbIGbrjN7gGxH4b8R+8FlhzbIJfvy1q637dFjRi9rJVmylRSOAB/fWPEzpx8zThmv
NqUJ3SP+EwI/H+5YzGCjJntU+dmzgXb0pVqKg8hwsDYxJHXPJAqR3SMI39VTC2uNBEV9vm57gGD1
9Z8anjesMJPNIY76J2fIBG3GVYA/yBsqRPgozmoqd9EF6DnaNoeVWTU098ZUaSTThZd+MUiXJs1Z
lT937Vb4wB05z5cTyD3OPcmQOnjlKodkGRG0aQXGl267QAt6UTEytXBjEACwoYl+iL56s1B9Ql98
Ne08gJHKqgKCfMxGL74c32p72iE43JKQrRR0MYz4izUC0vomASAm/AEt5IDYpK+0YiNpThmnoQ6t
JJqFeT2kys2RrPSjh+xTnTFrTSSeAPnSmLdgYmGS8ENtlhZcmhTA2EaASehlDJ/iPCCaTLKTQjyi
eUhzDueC/PNf8zF62kP2zSO47X97d0ZKmABFogJbRzlOgD4gLAZGizH9nRcMVna3GXxZ2Ns2y/+k
BRuHfI70lsOzRAfoNcb3Zk3v9cdf+Z0m8rjEWv8eIjI3bjEXCS7ZXAEyIxFSr2eg77v/JbYs3s0w
ssCi9iE31TmWf4VzlwFPJzH784AJtJW764LD7i3CRAdfCtLK22UR4772m6YlRYuCENxYgAe4OuMe
Axs70G7XJJZjahYKWR7elZOpfIFlJY4sqVp2/F71fVCbLarSD8EtEKyRY3CK2hpqQPA9x5UDZBMU
aFnqY/Yd2kDSZRO3KgD8pZSEUJx5v/lwGn07AFKDqhGa6ul4JknjDqM2z5Lr06/xFefHngk34UJt
nLWmWI9ALljeq5JaLvRWXf+ejghpd1+2/2pbggQJFqAw2V6Ujjv2ANCZG1tIhxVumb7DmVigTuv/
YuwuM4IW8mXdigmZyU2LZkmBU62fl3iKQToW2IgREf4yelGKNltcJy5f5tmmTsRYM5LbNar4X9yt
5dKtK3DWMPGE8y34l+kySIP6T3CccINoF5aQ2HMQ45S84lG3TnpzwUIHe+S1mvCGPV4Ymu3JvLhm
RIM1xpF9m9Rf
`pragma protect end_protected
