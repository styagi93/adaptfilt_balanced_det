��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR���[{�T���CK��TC,���:�
&��d!��]9�'D`�"9 S%�aQ�`!�6������V�W�l�a锦E(�\gC�slu�4U5=1�N�m��l�9ў��P���B�@+yg��=�}|��vFl�)TH�|/�gQ�T �����dn���l��IO���M�[n�K��y��=�'Nm���� �Tȓ�e�Da��"�1: ����);�5��`�y�0V<���1ڻϋ�h�=�H��Y�Lf��B���ce����+� ��~�kY�ա���lnT�V�dB!fw[t�|�I�t���1�'��)U�qE�zN�Ƌy5�jQ��r�ʷ�`⎬�lC@��TL㌠ ����f�� �`���ߛі����S���)
{H��
�ʑ����˂D�b�f�*���<R�>����{���ن���/2���T�[����V��K��mu���ڦF;��=�������F���i:�ّ��Yl7�V�%y3U!]O�8�$��n��j�6s+����^���s��$���@������/]C?)�g4�rxI����33"�'x*����PPy�d��8`�]�R�^VN�"��OCƕ(�'Υyl�դ��֩Q-(�ו�i9آ�l��4�7����&7�d��_yw'�"���'ü�����us0�d\}J#Q�4^L���E�Fy
1%O�6^j�A�M�����6�9�Ϥs�c�����ϒH�����R`��#��F���R�P�ę���qa����yu @`�'��H5�9䀙��0�e]
��;�� ?�4�X&�����<Z�/%�%���Np���>��O�:�nʅ��5��-�Յ)?�������Ht�s;
!��m�l�J��FY.�Ε����B��~b�N�9+�L&]z���|��w+�­H�5��Y'>ԗ��."$�����m\���k�)���f�]�TS���ϥ
;�Q���6zr	>*?��Ե�Jl���u �p�.O��d0��+w$#���L/�K�b��Y�X$��C?���F���{�2�jg�+�胃@���#-g�U���,�w8��ƕ�m~�	U����&U8{��-��������x㼱�N�JI)b&����nD��/��ZpJp���'/�+����[�!�1,e�y�4m�9�<�BLao~#��,�C�/��{�%V$�V����tZ�C8w}F̵�Mm�u�hk*�ٜ�.�\��(ÿ�K̀aɬ0C��9o�ю$4��_g񫺈)�F�|$�����K�\�v�]�@���vRh���-/��T�|'�3�3x�l(�"���rԃ�O��Ƨ-H�Ҁ���y0���W��/p���yh��+����N����%1����G;%��JLbAz�hۯ�z��7�ǚm���
.����@���f����t��H[��-U��>��+�����<F��bu�[�b����,�Ks�t�?�K��F�Y��� V�>,��(��u�k�±�a����?+"J�x���4xc��3Q\" �M�dO4$�V���
��F]hO��_mQt9�K{ZeD�͠�i1-�؛27aв�U3N���FR^zʁ�8C:Լf��>B>0�$�k*v択�ܙ$o��z8_0�:�,��Z���ޣ��SB�:�٬%7�I�F�s��Y`�eVw�qKp��d��)m����\XT���;¯ �^��#�&P��`S��7�B	s����L3�$�� ]���S|�9W���3�T^����smjA�g���>%�����Tc����/��z��Ǜ��{�w�sA|��������B<�3
`��~��؁��llվ�0�W*1b�#|��r�P_�k��B���5�e�A�y/D���}�&�Ml;�u����g�{Lu�|qE��J���;Y���Vl6�x�`�ܩ��x#tb�O�<�/ގ�W��PW8�(��gG� �Ӈ�>Ŝ-�|��fe���*���
���Q�q�h�>��h�)Zd��P�W��ࡐ(�eF(�HK;���Z����9�Z���a/�m%�E��k�en�:�:�ҥ9��>d �:@��e���{���о'z/��92�B1jX��e�Hd�2Mx�a��{�+���Fӿ��%�ttָ)$�T#�'�~�d�
�PãZK�V��W��(	��*p��� �BKk��38�jO.2��y10�e�_�\쨽C h�"C��`��bRH6� �_;�i7���� эl��˪>���H��t��g�?�mq�G���b�%*u ����'SV�$�gb�$7��T�o 0��h���U�]��5ß�Y�:&+q;�^��E�5O�3�'�x������R�ș�D�=ѿ'�(�2"�*Q�k(A�u� x��<S�K��7��NC��{B2W&�f V�W�G��W��v���r����ۈoy��(��q����(��RԻG�	��N1��T���<CE< qMfB����Je��S�!��'����<�`P�����������l��N���m���p^�D+$��OP���e��=��ݰ����9Z������Z+9�#����Au���5�"�����ׂ���Yv8��_��P�J̵�\i�A,[��g��9��k��D��OS�Ta��B�l�;�t� �GV��:5��K\G(5%e9����jP#�UV�x��@O����i�"�nàs��t9�_�g��U��Y×�o��[�Gt��+���\�?`�R�H-`\�Jִź҈/�nbz�#n����d��J�bw�(n,9c}��0?��e�!~�|�v���0�d���y�9��Hf�7���W|�ڈ4q��*{p4Y�g����%��o�U���ة?�]u#_lD=JZ�� U�SǑK��0[46GHۘo�<��>�察c�/���
ST6�'����H	�	�+�z������s
�̖y���9zY{V��� �S�63R��Lᄥ���$�	�� ����ӻm^��h�z�	�#���*���6hGK߄�#I�'�B�\���, �r��V�i�YuP`�L=��31����~��=�i�sqn�Y�8�����U��i��SO*"�}�?��|�h��7C�W�T���E!�S��N�r�4dV�啚=�gd�:
<F���c4��h�2
�/�O.���kẏ�So����\�!�]vpI��1�1�� �1��ËsZږ1eV��KZ22�aZs�G��6:øU9?��[Zt�4THLUh��ד����8'��d)=�J�)���8�h��X��:���T�=⊤��0N���䦛Nd��ݯ��ẃ�>�jA�F���4I�m��%���l$�ت5���Ψ���*�4m�"�8����,'v��P>L����om2X9,]o�����M82�o~�ד�@\��B�i�B��'8Y[D��LW��W�t��O�ڳú�m�lVJe�:B:�E��;o�����Wy��(T�s0� D�]II_�QK#�3�}�L/5���h�j�8;^�)�_��,@��
�gX~�7G ,)�ydq��r�I:w*%TX�D,�&b6ؠ}��c,V<LmwA��ed�h���/�%��F퍛��RHw�y����_mi#��V�uHd� �9Y�H�9,Pp��g}��V���T��~�0�9�у<��ޱ���e戀%���r6d�.n�~�	�d<�$�B*����U��	u��B uᕄg˭
!"r��Q����ĽX	 ��n�4��7b���rn�9{9:�b;�11Rh_��W,;����D�)�ʽ���_�O��E�ymeԊ-q�L�Z����C��>��)"����Mm�2�<�H�$-3����͹+Ϸ#&s�DQb g�� :��J�!� �:��v����нG��ഖU�Pk0r)Ī���hM��`�"Y�O�|&�ۿ��r��d86c�\FW�K�����"x6۬�2(_�	8.d��m�g���{,����sԱ�oW��S%�Ba��Y�R���uʅ�̶I3�3qa�/Sb�ӵ&%A��\�D�}�O�^�>U&��U/IY`�꒹�ν���i*�y���7@!�0&kQ��D��y �jT0%[{S2�Sn|6s8�Վb;-�7�!ƍ`�i�Z�ҹ ��^J�_�A1��b��4�ѳ�����{4����p��my���鉨�ut�6�Q�����b��K�˖L�l�	�ig��n� ˑ�bF���� -ళl��%,u8�I��аieqj�.�gRs)Ppy7�Pk�����h���c���֦)���ͿO���.7�)��ݛ��i4�@B��ȩ�ս{�x���Sn\X�Vp� �F1�UJ��xKv�W �0p��xW.v8Ea���.`�l� &�38��!���	B{"�0Wj}l�SRճ� �R>�(p�<:o��s�3m�����\
�N��u�H��N0=�|%�I�cG�AX�Jr#Б�;��c-��@�gN�a7u؂�wx+s���ￃ$=Z�!d#u0\ ����#�`U���͝��8���������1* [D�_���1eaX ��,?��z���yc�=�Y�?��R>����H'�]$�٥d�T�_�	��A�9o�0(�x��?�/p���,s�Y�Y�T �c���a|����p�'�@�>\f�p�<t�"���.�J�&=v�'�1��^�{��I1�KЏ�|�zR�;��B�	h��x_�8���1i!uB���0����� mB�	�Ό�г�ȒozK���9R"���%W��eY�JM[g@�F�[0Nq=�H��i��kQ{9��'�ʸ�+��0 �}hmUl$FM	S�Qjڂ���	0�2PJ�N��z:bݭ�Se�`Et�����rƳq�A>������]>)���^��,iu���Thd�~X)��j���^C��DU�+����w8٦[�>2��I��BЮ�#����^?m���ﱭo��Ŏ5ޚ`g�1��R�U|��W�Hf�A��6NWD�2��FT�%o~5(s�V@��qwW�[���x�t���j�#ԡc�X�2rc�<"�p���K?���;ڦb�`�`��?�M*?P��/���}�zĠ�B��i@�����P��l��hVŊS��l��a[���m�pH���D3L��ǥ��	�j��p���OY�в�5	ǟ�r��8�YMO�u:�U�F�n<��c��=jn'��a�7b_���X]�`��]%<�����d�5����9��3w�${�D�β��Z��j8_�R�U.ߍ���1a0�r�z&@�#��)�6_O��9βOGB�8~pR])(0A�qm�41�bN浍���o��wq`�kռ2���uҸEԐQ<���W�BNwl�i�xB`0V�͡�U'/�l���Q˲x��R ��;�b*]���V�����Jh��;�l?8��w�b����{�)%Uk�qu�{-�W��6�9k�9D����^�Ze��fNQ.��P��$�@/�O< �#���P~�5u]	����)�Ņ<Sx��u����CA[�9ZtV�'�[F��J�5 3�	d)��]pd�d�� `�~��Zۥ��p����@*Ψ)�ˀ�\��٦J���ݻHZ�ǐw����ĭ/�82��w19۞�����ráӍ�.����WJ�r�-5XP����;��1D���/oos���+����B�/��N�\���a���B���S{��W�����Eޫ�pN�1B\Qift	%�K�96��=w��T2(����]N0�FeJ�
!������f�Z0�%���_ux]�%�s����=e�m3��[2��Z�J��,��å��ͨ���?`����Y$J:����b��Z6&�3�}h�<��\a&[m��S���` ���*���I�+|Ẹ�/D���i�;�3 {�uU���.`)��|�5����Epe����5,�1~N��,ms>����\q́˒��������î�h�R[�a �'��*���nX��<-��X�����ף:�bu����e]��Zl\�٭�Y:,���B�}��)��Lj7Dɩz�n�e�Fh/<���Y���es�2=��Wg���l����e���x�[�] �nR�Ee;�\�ު��8����e�+��$�h�x����/6߱�&������߬^��ϫ�(�e/Jr7O�Ov�����L+4�)�\N�tp"�e?6������U ħ��hۤy��Q/���L7�W��0�~ĽQ�w\j�x���:	�+b����)�����G��0,��q z���,ߓ����õ Z��դ��t����]$#��6�bD�v'�k�K8͜�1ܳb�jx
�x��A��1���#��#ҿ�m%�;-�ԯ�P�8Ȩ��F0rv22���/�n{�]SpGn5apR�����&$+�QmI�a����4zOV��w_3,ư�����$���{�,_=(&���(���T�v;����ȣq���J�v��..J�X���DABit6����L�G ���H�)�Hq�wshl�#�4��=z��1��_��~qg%��i[ΦG=�._|"4��Ƙ���5�`�����`F���=v���Y�ն�gτy���P��V���m`]���%I�׳��4'afK�.,T�?	V����N�u*�ƶ��$S��7eShdͨ[v���`C�U��L	��:��}3<�u;���k[�?����k�\�u#�U��vXu9{��W����z,c�R����v�"��2�1qz
�-�K���h�Qyn������:B\��z��(�RD� ��}R�6 tK"Uq9v[��hv����$+�8