// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 16.0.0 Build 211 04/27/2016 SJ Lite Edition"

// DATE "04/14/2017 18:40:16"

// 
// Device: Altera EP4CE115F29C7 Package FBGA780
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module CIC (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	in_error,
	in_valid,
	in_ready,
	in0_data,
	in1_data,
	in2_data,
	in3_data,
	in4_data,
	in5_data,
	in6_data,
	in7_data,
	in8_data,
	in9_data,
	in10_data,
	in11_data,
	in12_data,
	in13_data,
	in14_data,
	in15_data,
	out_data,
	out_error,
	out_valid,
	out_ready,
	out_startofpacket,
	out_endofpacket,
	out_channel,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	[1:0] in_error;
input 	in_valid;
output 	in_ready;
input 	[15:0] in0_data;
input 	[15:0] in1_data;
input 	[15:0] in2_data;
input 	[15:0] in3_data;
input 	[15:0] in4_data;
input 	[15:0] in5_data;
input 	[15:0] in6_data;
input 	[15:0] in7_data;
input 	[15:0] in8_data;
input 	[15:0] in9_data;
input 	[15:0] in10_data;
input 	[15:0] in11_data;
input 	[15:0] in12_data;
input 	[15:0] in13_data;
input 	[15:0] in14_data;
input 	[15:0] in15_data;
output 	[15:0] out_data;
output 	[1:0] out_error;
output 	out_valid;
input 	out_ready;
output 	out_startofpacket;
output 	out_endofpacket;
output 	[3:0] out_channel;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \cic_ii_0|core|output_source_1|source_valid_s~q ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \cic_ii_0|out_data[0]~combout ;
wire \cic_ii_0|out_data[1]~combout ;
wire \cic_ii_0|out_data[2]~combout ;
wire \cic_ii_0|out_data[3]~combout ;
wire \cic_ii_0|out_data[4]~combout ;
wire \cic_ii_0|out_data[5]~combout ;
wire \cic_ii_0|out_data[6]~combout ;
wire \cic_ii_0|out_data[7]~combout ;
wire \cic_ii_0|out_data[8]~combout ;
wire \cic_ii_0|out_data[9]~combout ;
wire \cic_ii_0|out_data[10]~combout ;
wire \cic_ii_0|out_data[11]~combout ;
wire \cic_ii_0|out_data[12]~combout ;
wire \cic_ii_0|out_data[13]~combout ;
wire \cic_ii_0|out_data[14]~combout ;
wire \cic_ii_0|out_data[15]~combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \in0_data[0]~input_o ;
wire \in0_data[1]~input_o ;
wire \in0_data[2]~input_o ;
wire \in0_data[3]~input_o ;
wire \in1_data[0]~input_o ;
wire \in1_data[1]~input_o ;
wire \in1_data[2]~input_o ;
wire \in1_data[3]~input_o ;
wire \in2_data[0]~input_o ;
wire \in2_data[1]~input_o ;
wire \in2_data[2]~input_o ;
wire \in2_data[3]~input_o ;
wire \in3_data[0]~input_o ;
wire \in3_data[1]~input_o ;
wire \in3_data[2]~input_o ;
wire \in3_data[3]~input_o ;
wire \in4_data[0]~input_o ;
wire \in4_data[1]~input_o ;
wire \in4_data[2]~input_o ;
wire \in4_data[3]~input_o ;
wire \in5_data[0]~input_o ;
wire \in5_data[1]~input_o ;
wire \in5_data[2]~input_o ;
wire \in5_data[3]~input_o ;
wire \in6_data[0]~input_o ;
wire \in6_data[1]~input_o ;
wire \in6_data[2]~input_o ;
wire \in6_data[3]~input_o ;
wire \in7_data[0]~input_o ;
wire \in7_data[1]~input_o ;
wire \in7_data[2]~input_o ;
wire \in7_data[3]~input_o ;
wire \in8_data[0]~input_o ;
wire \in8_data[1]~input_o ;
wire \in8_data[2]~input_o ;
wire \in8_data[3]~input_o ;
wire \in9_data[0]~input_o ;
wire \in9_data[1]~input_o ;
wire \in9_data[2]~input_o ;
wire \in9_data[3]~input_o ;
wire \in10_data[0]~input_o ;
wire \in10_data[1]~input_o ;
wire \in10_data[2]~input_o ;
wire \in10_data[3]~input_o ;
wire \in11_data[0]~input_o ;
wire \in11_data[1]~input_o ;
wire \in11_data[2]~input_o ;
wire \in11_data[3]~input_o ;
wire \in12_data[0]~input_o ;
wire \in12_data[1]~input_o ;
wire \in12_data[2]~input_o ;
wire \in12_data[3]~input_o ;
wire \in13_data[0]~input_o ;
wire \in13_data[1]~input_o ;
wire \in13_data[2]~input_o ;
wire \in13_data[3]~input_o ;
wire \in14_data[0]~input_o ;
wire \in14_data[1]~input_o ;
wire \in14_data[2]~input_o ;
wire \in14_data[3]~input_o ;
wire \in15_data[0]~input_o ;
wire \in15_data[1]~input_o ;
wire \in15_data[2]~input_o ;
wire \in15_data[3]~input_o ;
wire \clk~input_o ;
wire \in_valid~input_o ;
wire \reset_n~input_o ;
wire \out_ready~input_o ;
wire \in10_data[10]~input_o ;
wire \in10_data[9]~input_o ;
wire \in10_data[8]~input_o ;
wire \in10_data[7]~input_o ;
wire \in10_data[6]~input_o ;
wire \in10_data[5]~input_o ;
wire \in10_data[4]~input_o ;
wire \in6_data[10]~input_o ;
wire \in6_data[9]~input_o ;
wire \in6_data[8]~input_o ;
wire \in6_data[7]~input_o ;
wire \in6_data[6]~input_o ;
wire \in6_data[5]~input_o ;
wire \in6_data[4]~input_o ;
wire \in14_data[10]~input_o ;
wire \in14_data[9]~input_o ;
wire \in14_data[8]~input_o ;
wire \in14_data[7]~input_o ;
wire \in14_data[6]~input_o ;
wire \in14_data[5]~input_o ;
wire \in14_data[4]~input_o ;
wire \in2_data[10]~input_o ;
wire \in2_data[9]~input_o ;
wire \in2_data[8]~input_o ;
wire \in2_data[7]~input_o ;
wire \in2_data[6]~input_o ;
wire \in2_data[5]~input_o ;
wire \in2_data[4]~input_o ;
wire \in11_data[10]~input_o ;
wire \in11_data[9]~input_o ;
wire \in11_data[8]~input_o ;
wire \in11_data[7]~input_o ;
wire \in11_data[6]~input_o ;
wire \in11_data[5]~input_o ;
wire \in11_data[4]~input_o ;
wire \in7_data[10]~input_o ;
wire \in7_data[9]~input_o ;
wire \in7_data[8]~input_o ;
wire \in7_data[7]~input_o ;
wire \in7_data[6]~input_o ;
wire \in7_data[5]~input_o ;
wire \in7_data[4]~input_o ;
wire \in15_data[10]~input_o ;
wire \in15_data[9]~input_o ;
wire \in15_data[8]~input_o ;
wire \in15_data[7]~input_o ;
wire \in15_data[6]~input_o ;
wire \in15_data[5]~input_o ;
wire \in15_data[4]~input_o ;
wire \in3_data[10]~input_o ;
wire \in3_data[9]~input_o ;
wire \in3_data[8]~input_o ;
wire \in3_data[7]~input_o ;
wire \in3_data[6]~input_o ;
wire \in3_data[5]~input_o ;
wire \in3_data[4]~input_o ;
wire \in5_data[10]~input_o ;
wire \in5_data[9]~input_o ;
wire \in5_data[8]~input_o ;
wire \in5_data[7]~input_o ;
wire \in5_data[6]~input_o ;
wire \in5_data[5]~input_o ;
wire \in5_data[4]~input_o ;
wire \in9_data[10]~input_o ;
wire \in9_data[9]~input_o ;
wire \in9_data[8]~input_o ;
wire \in9_data[7]~input_o ;
wire \in9_data[6]~input_o ;
wire \in9_data[5]~input_o ;
wire \in9_data[4]~input_o ;
wire \in13_data[10]~input_o ;
wire \in13_data[9]~input_o ;
wire \in13_data[8]~input_o ;
wire \in13_data[7]~input_o ;
wire \in13_data[6]~input_o ;
wire \in13_data[5]~input_o ;
wire \in13_data[4]~input_o ;
wire \in1_data[10]~input_o ;
wire \in1_data[9]~input_o ;
wire \in1_data[8]~input_o ;
wire \in1_data[7]~input_o ;
wire \in1_data[6]~input_o ;
wire \in1_data[5]~input_o ;
wire \in1_data[4]~input_o ;
wire \in4_data[10]~input_o ;
wire \in4_data[9]~input_o ;
wire \in4_data[8]~input_o ;
wire \in4_data[7]~input_o ;
wire \in4_data[6]~input_o ;
wire \in4_data[5]~input_o ;
wire \in4_data[4]~input_o ;
wire \in8_data[10]~input_o ;
wire \in8_data[9]~input_o ;
wire \in8_data[8]~input_o ;
wire \in8_data[7]~input_o ;
wire \in8_data[6]~input_o ;
wire \in8_data[5]~input_o ;
wire \in8_data[4]~input_o ;
wire \in12_data[10]~input_o ;
wire \in12_data[9]~input_o ;
wire \in12_data[8]~input_o ;
wire \in12_data[7]~input_o ;
wire \in12_data[6]~input_o ;
wire \in12_data[5]~input_o ;
wire \in12_data[4]~input_o ;
wire \in0_data[10]~input_o ;
wire \in0_data[9]~input_o ;
wire \in0_data[8]~input_o ;
wire \in0_data[7]~input_o ;
wire \in0_data[6]~input_o ;
wire \in0_data[5]~input_o ;
wire \in0_data[4]~input_o ;
wire \in6_data[11]~input_o ;
wire \in7_data[11]~input_o ;
wire \in5_data[11]~input_o ;
wire \in4_data[11]~input_o ;
wire \in10_data[11]~input_o ;
wire \in11_data[11]~input_o ;
wire \in9_data[11]~input_o ;
wire \in8_data[11]~input_o ;
wire \in14_data[11]~input_o ;
wire \in15_data[11]~input_o ;
wire \in13_data[11]~input_o ;
wire \in12_data[11]~input_o ;
wire \in2_data[11]~input_o ;
wire \in3_data[11]~input_o ;
wire \in1_data[11]~input_o ;
wire \in0_data[11]~input_o ;
wire \in6_data[12]~input_o ;
wire \in10_data[12]~input_o ;
wire \in14_data[12]~input_o ;
wire \in2_data[12]~input_o ;
wire \in7_data[12]~input_o ;
wire \in11_data[12]~input_o ;
wire \in15_data[12]~input_o ;
wire \in3_data[12]~input_o ;
wire \in9_data[12]~input_o ;
wire \in5_data[12]~input_o ;
wire \in13_data[12]~input_o ;
wire \in1_data[12]~input_o ;
wire \in8_data[12]~input_o ;
wire \in4_data[12]~input_o ;
wire \in12_data[12]~input_o ;
wire \in0_data[12]~input_o ;
wire \in10_data[13]~input_o ;
wire \in11_data[13]~input_o ;
wire \in9_data[13]~input_o ;
wire \in8_data[13]~input_o ;
wire \in6_data[13]~input_o ;
wire \in7_data[13]~input_o ;
wire \in5_data[13]~input_o ;
wire \in4_data[13]~input_o ;
wire \in14_data[13]~input_o ;
wire \in15_data[13]~input_o ;
wire \in13_data[13]~input_o ;
wire \in12_data[13]~input_o ;
wire \in2_data[13]~input_o ;
wire \in3_data[13]~input_o ;
wire \in1_data[13]~input_o ;
wire \in0_data[13]~input_o ;
wire \in10_data[14]~input_o ;
wire \in6_data[14]~input_o ;
wire \in14_data[14]~input_o ;
wire \in2_data[14]~input_o ;
wire \in11_data[14]~input_o ;
wire \in7_data[14]~input_o ;
wire \in15_data[14]~input_o ;
wire \in3_data[14]~input_o ;
wire \in5_data[14]~input_o ;
wire \in9_data[14]~input_o ;
wire \in13_data[14]~input_o ;
wire \in1_data[14]~input_o ;
wire \in4_data[14]~input_o ;
wire \in8_data[14]~input_o ;
wire \in12_data[14]~input_o ;
wire \in0_data[14]~input_o ;
wire \in6_data[15]~input_o ;
wire \in7_data[15]~input_o ;
wire \in5_data[15]~input_o ;
wire \in4_data[15]~input_o ;
wire \in10_data[15]~input_o ;
wire \in11_data[15]~input_o ;
wire \in9_data[15]~input_o ;
wire \in8_data[15]~input_o ;
wire \in14_data[15]~input_o ;
wire \in15_data[15]~input_o ;
wire \in13_data[15]~input_o ;
wire \in12_data[15]~input_o ;
wire \in2_data[15]~input_o ;
wire \in3_data[15]~input_o ;
wire \in1_data[15]~input_o ;
wire \in0_data[15]~input_o ;
wire \in_error[0]~input_o ;
wire \in_error[1]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \~GND~combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~1 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~3 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~5 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~7 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~3_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


CIC_CIC_cic_ii_0 cic_ii_0(
	.full_dff(\cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ),
	.source_valid_s(\cic_ii_0|core|output_source_1|source_valid_s~q ),
	.q_b_16(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_17(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_18(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_19(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.out_data_0(\cic_ii_0|out_data[0]~combout ),
	.out_data_1(\cic_ii_0|out_data[1]~combout ),
	.out_data_2(\cic_ii_0|out_data[2]~combout ),
	.out_data_3(\cic_ii_0|out_data[3]~combout ),
	.out_data_4(\cic_ii_0|out_data[4]~combout ),
	.out_data_5(\cic_ii_0|out_data[5]~combout ),
	.out_data_6(\cic_ii_0|out_data[6]~combout ),
	.out_data_7(\cic_ii_0|out_data[7]~combout ),
	.out_data_8(\cic_ii_0|out_data[8]~combout ),
	.out_data_9(\cic_ii_0|out_data[9]~combout ),
	.out_data_10(\cic_ii_0|out_data[10]~combout ),
	.out_data_11(\cic_ii_0|out_data[11]~combout ),
	.out_data_12(\cic_ii_0|out_data[12]~combout ),
	.out_data_13(\cic_ii_0|out_data[13]~combout ),
	.out_data_14(\cic_ii_0|out_data[14]~combout ),
	.out_data_15(\cic_ii_0|out_data[15]~combout ),
	.GND_port(\~GND~combout ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.clk(\clk~input_o ),
	.in_valid(\in_valid~input_o ),
	.reset_n(\reset_n~input_o ),
	.out_ready(\out_ready~input_o ),
	.in10_data_10(\in10_data[10]~input_o ),
	.in10_data_9(\in10_data[9]~input_o ),
	.in10_data_8(\in10_data[8]~input_o ),
	.in10_data_7(\in10_data[7]~input_o ),
	.in10_data_6(\in10_data[6]~input_o ),
	.in10_data_5(\in10_data[5]~input_o ),
	.in10_data_4(\in10_data[4]~input_o ),
	.in6_data_10(\in6_data[10]~input_o ),
	.in6_data_9(\in6_data[9]~input_o ),
	.in6_data_8(\in6_data[8]~input_o ),
	.in6_data_7(\in6_data[7]~input_o ),
	.in6_data_6(\in6_data[6]~input_o ),
	.in6_data_5(\in6_data[5]~input_o ),
	.in6_data_4(\in6_data[4]~input_o ),
	.in14_data_10(\in14_data[10]~input_o ),
	.in14_data_9(\in14_data[9]~input_o ),
	.in14_data_8(\in14_data[8]~input_o ),
	.in14_data_7(\in14_data[7]~input_o ),
	.in14_data_6(\in14_data[6]~input_o ),
	.in14_data_5(\in14_data[5]~input_o ),
	.in14_data_4(\in14_data[4]~input_o ),
	.in2_data_10(\in2_data[10]~input_o ),
	.in2_data_9(\in2_data[9]~input_o ),
	.in2_data_8(\in2_data[8]~input_o ),
	.in2_data_7(\in2_data[7]~input_o ),
	.in2_data_6(\in2_data[6]~input_o ),
	.in2_data_5(\in2_data[5]~input_o ),
	.in2_data_4(\in2_data[4]~input_o ),
	.in11_data_10(\in11_data[10]~input_o ),
	.in11_data_9(\in11_data[9]~input_o ),
	.in11_data_8(\in11_data[8]~input_o ),
	.in11_data_7(\in11_data[7]~input_o ),
	.in11_data_6(\in11_data[6]~input_o ),
	.in11_data_5(\in11_data[5]~input_o ),
	.in11_data_4(\in11_data[4]~input_o ),
	.in7_data_10(\in7_data[10]~input_o ),
	.in7_data_9(\in7_data[9]~input_o ),
	.in7_data_8(\in7_data[8]~input_o ),
	.in7_data_7(\in7_data[7]~input_o ),
	.in7_data_6(\in7_data[6]~input_o ),
	.in7_data_5(\in7_data[5]~input_o ),
	.in7_data_4(\in7_data[4]~input_o ),
	.in15_data_10(\in15_data[10]~input_o ),
	.in15_data_9(\in15_data[9]~input_o ),
	.in15_data_8(\in15_data[8]~input_o ),
	.in15_data_7(\in15_data[7]~input_o ),
	.in15_data_6(\in15_data[6]~input_o ),
	.in15_data_5(\in15_data[5]~input_o ),
	.in15_data_4(\in15_data[4]~input_o ),
	.in3_data_10(\in3_data[10]~input_o ),
	.in3_data_9(\in3_data[9]~input_o ),
	.in3_data_8(\in3_data[8]~input_o ),
	.in3_data_7(\in3_data[7]~input_o ),
	.in3_data_6(\in3_data[6]~input_o ),
	.in3_data_5(\in3_data[5]~input_o ),
	.in3_data_4(\in3_data[4]~input_o ),
	.in5_data_10(\in5_data[10]~input_o ),
	.in5_data_9(\in5_data[9]~input_o ),
	.in5_data_8(\in5_data[8]~input_o ),
	.in5_data_7(\in5_data[7]~input_o ),
	.in5_data_6(\in5_data[6]~input_o ),
	.in5_data_5(\in5_data[5]~input_o ),
	.in5_data_4(\in5_data[4]~input_o ),
	.in9_data_10(\in9_data[10]~input_o ),
	.in9_data_9(\in9_data[9]~input_o ),
	.in9_data_8(\in9_data[8]~input_o ),
	.in9_data_7(\in9_data[7]~input_o ),
	.in9_data_6(\in9_data[6]~input_o ),
	.in9_data_5(\in9_data[5]~input_o ),
	.in9_data_4(\in9_data[4]~input_o ),
	.in13_data_10(\in13_data[10]~input_o ),
	.in13_data_9(\in13_data[9]~input_o ),
	.in13_data_8(\in13_data[8]~input_o ),
	.in13_data_7(\in13_data[7]~input_o ),
	.in13_data_6(\in13_data[6]~input_o ),
	.in13_data_5(\in13_data[5]~input_o ),
	.in13_data_4(\in13_data[4]~input_o ),
	.in1_data_10(\in1_data[10]~input_o ),
	.in1_data_9(\in1_data[9]~input_o ),
	.in1_data_8(\in1_data[8]~input_o ),
	.in1_data_7(\in1_data[7]~input_o ),
	.in1_data_6(\in1_data[6]~input_o ),
	.in1_data_5(\in1_data[5]~input_o ),
	.in1_data_4(\in1_data[4]~input_o ),
	.in4_data_10(\in4_data[10]~input_o ),
	.in4_data_9(\in4_data[9]~input_o ),
	.in4_data_8(\in4_data[8]~input_o ),
	.in4_data_7(\in4_data[7]~input_o ),
	.in4_data_6(\in4_data[6]~input_o ),
	.in4_data_5(\in4_data[5]~input_o ),
	.in4_data_4(\in4_data[4]~input_o ),
	.in8_data_10(\in8_data[10]~input_o ),
	.in8_data_9(\in8_data[9]~input_o ),
	.in8_data_8(\in8_data[8]~input_o ),
	.in8_data_7(\in8_data[7]~input_o ),
	.in8_data_6(\in8_data[6]~input_o ),
	.in8_data_5(\in8_data[5]~input_o ),
	.in8_data_4(\in8_data[4]~input_o ),
	.in12_data_10(\in12_data[10]~input_o ),
	.in12_data_9(\in12_data[9]~input_o ),
	.in12_data_8(\in12_data[8]~input_o ),
	.in12_data_7(\in12_data[7]~input_o ),
	.in12_data_6(\in12_data[6]~input_o ),
	.in12_data_5(\in12_data[5]~input_o ),
	.in12_data_4(\in12_data[4]~input_o ),
	.in0_data_10(\in0_data[10]~input_o ),
	.in0_data_9(\in0_data[9]~input_o ),
	.in0_data_8(\in0_data[8]~input_o ),
	.in0_data_7(\in0_data[7]~input_o ),
	.in0_data_6(\in0_data[6]~input_o ),
	.in0_data_5(\in0_data[5]~input_o ),
	.in0_data_4(\in0_data[4]~input_o ),
	.in6_data_11(\in6_data[11]~input_o ),
	.in7_data_11(\in7_data[11]~input_o ),
	.in5_data_11(\in5_data[11]~input_o ),
	.in4_data_11(\in4_data[11]~input_o ),
	.in10_data_11(\in10_data[11]~input_o ),
	.in11_data_11(\in11_data[11]~input_o ),
	.in9_data_11(\in9_data[11]~input_o ),
	.in8_data_11(\in8_data[11]~input_o ),
	.in14_data_11(\in14_data[11]~input_o ),
	.in15_data_11(\in15_data[11]~input_o ),
	.in13_data_11(\in13_data[11]~input_o ),
	.in12_data_11(\in12_data[11]~input_o ),
	.in2_data_11(\in2_data[11]~input_o ),
	.in3_data_11(\in3_data[11]~input_o ),
	.in1_data_11(\in1_data[11]~input_o ),
	.in0_data_11(\in0_data[11]~input_o ),
	.in6_data_12(\in6_data[12]~input_o ),
	.in10_data_12(\in10_data[12]~input_o ),
	.in14_data_12(\in14_data[12]~input_o ),
	.in2_data_12(\in2_data[12]~input_o ),
	.in7_data_12(\in7_data[12]~input_o ),
	.in11_data_12(\in11_data[12]~input_o ),
	.in15_data_12(\in15_data[12]~input_o ),
	.in3_data_12(\in3_data[12]~input_o ),
	.in9_data_12(\in9_data[12]~input_o ),
	.in5_data_12(\in5_data[12]~input_o ),
	.in13_data_12(\in13_data[12]~input_o ),
	.in1_data_12(\in1_data[12]~input_o ),
	.in8_data_12(\in8_data[12]~input_o ),
	.in4_data_12(\in4_data[12]~input_o ),
	.in12_data_12(\in12_data[12]~input_o ),
	.in0_data_12(\in0_data[12]~input_o ),
	.in10_data_13(\in10_data[13]~input_o ),
	.in11_data_13(\in11_data[13]~input_o ),
	.in9_data_13(\in9_data[13]~input_o ),
	.in8_data_13(\in8_data[13]~input_o ),
	.in6_data_13(\in6_data[13]~input_o ),
	.in7_data_13(\in7_data[13]~input_o ),
	.in5_data_13(\in5_data[13]~input_o ),
	.in4_data_13(\in4_data[13]~input_o ),
	.in14_data_13(\in14_data[13]~input_o ),
	.in15_data_13(\in15_data[13]~input_o ),
	.in13_data_13(\in13_data[13]~input_o ),
	.in12_data_13(\in12_data[13]~input_o ),
	.in2_data_13(\in2_data[13]~input_o ),
	.in3_data_13(\in3_data[13]~input_o ),
	.in1_data_13(\in1_data[13]~input_o ),
	.in0_data_13(\in0_data[13]~input_o ),
	.in10_data_14(\in10_data[14]~input_o ),
	.in6_data_14(\in6_data[14]~input_o ),
	.in14_data_14(\in14_data[14]~input_o ),
	.in2_data_14(\in2_data[14]~input_o ),
	.in11_data_14(\in11_data[14]~input_o ),
	.in7_data_14(\in7_data[14]~input_o ),
	.in15_data_14(\in15_data[14]~input_o ),
	.in3_data_14(\in3_data[14]~input_o ),
	.in5_data_14(\in5_data[14]~input_o ),
	.in9_data_14(\in9_data[14]~input_o ),
	.in13_data_14(\in13_data[14]~input_o ),
	.in1_data_14(\in1_data[14]~input_o ),
	.in4_data_14(\in4_data[14]~input_o ),
	.in8_data_14(\in8_data[14]~input_o ),
	.in12_data_14(\in12_data[14]~input_o ),
	.in0_data_14(\in0_data[14]~input_o ),
	.in6_data_15(\in6_data[15]~input_o ),
	.in7_data_15(\in7_data[15]~input_o ),
	.in5_data_15(\in5_data[15]~input_o ),
	.in4_data_15(\in4_data[15]~input_o ),
	.in10_data_15(\in10_data[15]~input_o ),
	.in11_data_15(\in11_data[15]~input_o ),
	.in9_data_15(\in9_data[15]~input_o ),
	.in8_data_15(\in8_data[15]~input_o ),
	.in14_data_15(\in14_data[15]~input_o ),
	.in15_data_15(\in15_data[15]~input_o ),
	.in13_data_15(\in13_data[15]~input_o ),
	.in12_data_15(\in12_data[15]~input_o ),
	.in2_data_15(\in2_data[15]~input_o ),
	.in3_data_15(\in3_data[15]~input_o ),
	.in1_data_15(\in1_data[15]~input_o ),
	.in0_data_15(\in0_data[15]~input_o ));

assign \clk~input_o  = clk;

assign \in_valid~input_o  = in_valid;

assign \reset_n~input_o  = reset_n;

assign \out_ready~input_o  = out_ready;

assign \in10_data[10]~input_o  = in10_data[10];

assign \in10_data[9]~input_o  = in10_data[9];

assign \in10_data[8]~input_o  = in10_data[8];

assign \in10_data[7]~input_o  = in10_data[7];

assign \in10_data[6]~input_o  = in10_data[6];

assign \in10_data[5]~input_o  = in10_data[5];

assign \in10_data[4]~input_o  = in10_data[4];

assign \in6_data[10]~input_o  = in6_data[10];

assign \in6_data[9]~input_o  = in6_data[9];

assign \in6_data[8]~input_o  = in6_data[8];

assign \in6_data[7]~input_o  = in6_data[7];

assign \in6_data[6]~input_o  = in6_data[6];

assign \in6_data[5]~input_o  = in6_data[5];

assign \in6_data[4]~input_o  = in6_data[4];

assign \in14_data[10]~input_o  = in14_data[10];

assign \in14_data[9]~input_o  = in14_data[9];

assign \in14_data[8]~input_o  = in14_data[8];

assign \in14_data[7]~input_o  = in14_data[7];

assign \in14_data[6]~input_o  = in14_data[6];

assign \in14_data[5]~input_o  = in14_data[5];

assign \in14_data[4]~input_o  = in14_data[4];

assign \in2_data[10]~input_o  = in2_data[10];

assign \in2_data[9]~input_o  = in2_data[9];

assign \in2_data[8]~input_o  = in2_data[8];

assign \in2_data[7]~input_o  = in2_data[7];

assign \in2_data[6]~input_o  = in2_data[6];

assign \in2_data[5]~input_o  = in2_data[5];

assign \in2_data[4]~input_o  = in2_data[4];

assign \in11_data[10]~input_o  = in11_data[10];

assign \in11_data[9]~input_o  = in11_data[9];

assign \in11_data[8]~input_o  = in11_data[8];

assign \in11_data[7]~input_o  = in11_data[7];

assign \in11_data[6]~input_o  = in11_data[6];

assign \in11_data[5]~input_o  = in11_data[5];

assign \in11_data[4]~input_o  = in11_data[4];

assign \in7_data[10]~input_o  = in7_data[10];

assign \in7_data[9]~input_o  = in7_data[9];

assign \in7_data[8]~input_o  = in7_data[8];

assign \in7_data[7]~input_o  = in7_data[7];

assign \in7_data[6]~input_o  = in7_data[6];

assign \in7_data[5]~input_o  = in7_data[5];

assign \in7_data[4]~input_o  = in7_data[4];

assign \in15_data[10]~input_o  = in15_data[10];

assign \in15_data[9]~input_o  = in15_data[9];

assign \in15_data[8]~input_o  = in15_data[8];

assign \in15_data[7]~input_o  = in15_data[7];

assign \in15_data[6]~input_o  = in15_data[6];

assign \in15_data[5]~input_o  = in15_data[5];

assign \in15_data[4]~input_o  = in15_data[4];

assign \in3_data[10]~input_o  = in3_data[10];

assign \in3_data[9]~input_o  = in3_data[9];

assign \in3_data[8]~input_o  = in3_data[8];

assign \in3_data[7]~input_o  = in3_data[7];

assign \in3_data[6]~input_o  = in3_data[6];

assign \in3_data[5]~input_o  = in3_data[5];

assign \in3_data[4]~input_o  = in3_data[4];

assign \in5_data[10]~input_o  = in5_data[10];

assign \in5_data[9]~input_o  = in5_data[9];

assign \in5_data[8]~input_o  = in5_data[8];

assign \in5_data[7]~input_o  = in5_data[7];

assign \in5_data[6]~input_o  = in5_data[6];

assign \in5_data[5]~input_o  = in5_data[5];

assign \in5_data[4]~input_o  = in5_data[4];

assign \in9_data[10]~input_o  = in9_data[10];

assign \in9_data[9]~input_o  = in9_data[9];

assign \in9_data[8]~input_o  = in9_data[8];

assign \in9_data[7]~input_o  = in9_data[7];

assign \in9_data[6]~input_o  = in9_data[6];

assign \in9_data[5]~input_o  = in9_data[5];

assign \in9_data[4]~input_o  = in9_data[4];

assign \in13_data[10]~input_o  = in13_data[10];

assign \in13_data[9]~input_o  = in13_data[9];

assign \in13_data[8]~input_o  = in13_data[8];

assign \in13_data[7]~input_o  = in13_data[7];

assign \in13_data[6]~input_o  = in13_data[6];

assign \in13_data[5]~input_o  = in13_data[5];

assign \in13_data[4]~input_o  = in13_data[4];

assign \in1_data[10]~input_o  = in1_data[10];

assign \in1_data[9]~input_o  = in1_data[9];

assign \in1_data[8]~input_o  = in1_data[8];

assign \in1_data[7]~input_o  = in1_data[7];

assign \in1_data[6]~input_o  = in1_data[6];

assign \in1_data[5]~input_o  = in1_data[5];

assign \in1_data[4]~input_o  = in1_data[4];

assign \in4_data[10]~input_o  = in4_data[10];

assign \in4_data[9]~input_o  = in4_data[9];

assign \in4_data[8]~input_o  = in4_data[8];

assign \in4_data[7]~input_o  = in4_data[7];

assign \in4_data[6]~input_o  = in4_data[6];

assign \in4_data[5]~input_o  = in4_data[5];

assign \in4_data[4]~input_o  = in4_data[4];

assign \in8_data[10]~input_o  = in8_data[10];

assign \in8_data[9]~input_o  = in8_data[9];

assign \in8_data[8]~input_o  = in8_data[8];

assign \in8_data[7]~input_o  = in8_data[7];

assign \in8_data[6]~input_o  = in8_data[6];

assign \in8_data[5]~input_o  = in8_data[5];

assign \in8_data[4]~input_o  = in8_data[4];

assign \in12_data[10]~input_o  = in12_data[10];

assign \in12_data[9]~input_o  = in12_data[9];

assign \in12_data[8]~input_o  = in12_data[8];

assign \in12_data[7]~input_o  = in12_data[7];

assign \in12_data[6]~input_o  = in12_data[6];

assign \in12_data[5]~input_o  = in12_data[5];

assign \in12_data[4]~input_o  = in12_data[4];

assign \in0_data[10]~input_o  = in0_data[10];

assign \in0_data[9]~input_o  = in0_data[9];

assign \in0_data[8]~input_o  = in0_data[8];

assign \in0_data[7]~input_o  = in0_data[7];

assign \in0_data[6]~input_o  = in0_data[6];

assign \in0_data[5]~input_o  = in0_data[5];

assign \in0_data[4]~input_o  = in0_data[4];

assign \in6_data[11]~input_o  = in6_data[11];

assign \in7_data[11]~input_o  = in7_data[11];

assign \in5_data[11]~input_o  = in5_data[11];

assign \in4_data[11]~input_o  = in4_data[11];

assign \in10_data[11]~input_o  = in10_data[11];

assign \in11_data[11]~input_o  = in11_data[11];

assign \in9_data[11]~input_o  = in9_data[11];

assign \in8_data[11]~input_o  = in8_data[11];

assign \in14_data[11]~input_o  = in14_data[11];

assign \in15_data[11]~input_o  = in15_data[11];

assign \in13_data[11]~input_o  = in13_data[11];

assign \in12_data[11]~input_o  = in12_data[11];

assign \in2_data[11]~input_o  = in2_data[11];

assign \in3_data[11]~input_o  = in3_data[11];

assign \in1_data[11]~input_o  = in1_data[11];

assign \in0_data[11]~input_o  = in0_data[11];

assign \in6_data[12]~input_o  = in6_data[12];

assign \in10_data[12]~input_o  = in10_data[12];

assign \in14_data[12]~input_o  = in14_data[12];

assign \in2_data[12]~input_o  = in2_data[12];

assign \in7_data[12]~input_o  = in7_data[12];

assign \in11_data[12]~input_o  = in11_data[12];

assign \in15_data[12]~input_o  = in15_data[12];

assign \in3_data[12]~input_o  = in3_data[12];

assign \in9_data[12]~input_o  = in9_data[12];

assign \in5_data[12]~input_o  = in5_data[12];

assign \in13_data[12]~input_o  = in13_data[12];

assign \in1_data[12]~input_o  = in1_data[12];

assign \in8_data[12]~input_o  = in8_data[12];

assign \in4_data[12]~input_o  = in4_data[12];

assign \in12_data[12]~input_o  = in12_data[12];

assign \in0_data[12]~input_o  = in0_data[12];

assign \in10_data[13]~input_o  = in10_data[13];

assign \in11_data[13]~input_o  = in11_data[13];

assign \in9_data[13]~input_o  = in9_data[13];

assign \in8_data[13]~input_o  = in8_data[13];

assign \in6_data[13]~input_o  = in6_data[13];

assign \in7_data[13]~input_o  = in7_data[13];

assign \in5_data[13]~input_o  = in5_data[13];

assign \in4_data[13]~input_o  = in4_data[13];

assign \in14_data[13]~input_o  = in14_data[13];

assign \in15_data[13]~input_o  = in15_data[13];

assign \in13_data[13]~input_o  = in13_data[13];

assign \in12_data[13]~input_o  = in12_data[13];

assign \in2_data[13]~input_o  = in2_data[13];

assign \in3_data[13]~input_o  = in3_data[13];

assign \in1_data[13]~input_o  = in1_data[13];

assign \in0_data[13]~input_o  = in0_data[13];

assign \in10_data[14]~input_o  = in10_data[14];

assign \in6_data[14]~input_o  = in6_data[14];

assign \in14_data[14]~input_o  = in14_data[14];

assign \in2_data[14]~input_o  = in2_data[14];

assign \in11_data[14]~input_o  = in11_data[14];

assign \in7_data[14]~input_o  = in7_data[14];

assign \in15_data[14]~input_o  = in15_data[14];

assign \in3_data[14]~input_o  = in3_data[14];

assign \in5_data[14]~input_o  = in5_data[14];

assign \in9_data[14]~input_o  = in9_data[14];

assign \in13_data[14]~input_o  = in13_data[14];

assign \in1_data[14]~input_o  = in1_data[14];

assign \in4_data[14]~input_o  = in4_data[14];

assign \in8_data[14]~input_o  = in8_data[14];

assign \in12_data[14]~input_o  = in12_data[14];

assign \in0_data[14]~input_o  = in0_data[14];

assign \in6_data[15]~input_o  = in6_data[15];

assign \in7_data[15]~input_o  = in7_data[15];

assign \in5_data[15]~input_o  = in5_data[15];

assign \in4_data[15]~input_o  = in4_data[15];

assign \in10_data[15]~input_o  = in10_data[15];

assign \in11_data[15]~input_o  = in11_data[15];

assign \in9_data[15]~input_o  = in9_data[15];

assign \in8_data[15]~input_o  = in8_data[15];

assign \in14_data[15]~input_o  = in14_data[15];

assign \in15_data[15]~input_o  = in15_data[15];

assign \in13_data[15]~input_o  = in13_data[15];

assign \in12_data[15]~input_o  = in12_data[15];

assign \in2_data[15]~input_o  = in2_data[15];

assign \in3_data[15]~input_o  = in3_data[15];

assign \in1_data[15]~input_o  = in1_data[15];

assign \in0_data[15]~input_o  = in0_data[15];

assign in_ready = ~ \cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ;

assign out_data[0] = \cic_ii_0|out_data[0]~combout ;

assign out_data[1] = \cic_ii_0|out_data[1]~combout ;

assign out_data[2] = \cic_ii_0|out_data[2]~combout ;

assign out_data[3] = \cic_ii_0|out_data[3]~combout ;

assign out_data[4] = \cic_ii_0|out_data[4]~combout ;

assign out_data[5] = \cic_ii_0|out_data[5]~combout ;

assign out_data[6] = \cic_ii_0|out_data[6]~combout ;

assign out_data[7] = \cic_ii_0|out_data[7]~combout ;

assign out_data[8] = \cic_ii_0|out_data[8]~combout ;

assign out_data[9] = \cic_ii_0|out_data[9]~combout ;

assign out_data[10] = \cic_ii_0|out_data[10]~combout ;

assign out_data[11] = \cic_ii_0|out_data[11]~combout ;

assign out_data[12] = \cic_ii_0|out_data[12]~combout ;

assign out_data[13] = \cic_ii_0|out_data[13]~combout ;

assign out_data[14] = \cic_ii_0|out_data[14]~combout ;

assign out_data[15] = \cic_ii_0|out_data[15]~combout ;

assign out_error[0] = \in_error[0]~input_o ;

assign out_error[1] = \in_error[1]~input_o ;

assign out_valid = \cic_ii_0|core|output_source_1|source_valid_s~q ;

assign out_startofpacket = gnd;

assign out_endofpacket = gnd;

assign out_channel[0] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;

assign out_channel[1] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;

assign out_channel[2] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;

assign out_channel[3] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \in_error[0]~input_o  = in_error[0];

assign \in_error[1]~input_o  = in_error[1];

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cycloneive_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 (
	.dataa(\~GND~combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .lut_mask = 16'hFEFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .lut_mask = 16'h7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3 .lut_mask = 16'hFEFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_1 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_2 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 16'hFDFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|AMGP4450~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|AMGP4450 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.datad(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~13 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'h6FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 16'hD8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .lut_mask = 16'h8BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .lut_mask = 16'h96FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~1 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0 .lut_mask = 16'h55AA;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 .lut_mask = 16'h9966;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~1 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~3 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2 .lut_mask = 16'h5A5F;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .lut_mask = 16'h9966;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~3 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~5 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4 .lut_mask = 16'h5AAF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4 .sum_lutc_input = "cin";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~5 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~7 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6 .lut_mask = 16'h5A5F;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6 .sum_lutc_input = "cin";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~7 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8 .lut_mask = 16'h5A5A;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .lut_mask = 16'h9966;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~0 .lut_mask = 16'hCC55;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5 .lut_mask = 16'hF6F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6 .lut_mask = 16'h66FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~1 .lut_mask = 16'hAACC;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~2 .lut_mask = 16'hAACC;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .lut_mask = 16'hF6FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~3 .lut_mask = 16'hAA33;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~2_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~1_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~0_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .sum_lutc_input = "datac";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

cycloneive_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|tdo~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

cycloneive_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

assign \in0_data[0]~input_o  = in0_data[0];

assign \in0_data[1]~input_o  = in0_data[1];

assign \in0_data[2]~input_o  = in0_data[2];

assign \in0_data[3]~input_o  = in0_data[3];

assign \in1_data[0]~input_o  = in1_data[0];

assign \in1_data[1]~input_o  = in1_data[1];

assign \in1_data[2]~input_o  = in1_data[2];

assign \in1_data[3]~input_o  = in1_data[3];

assign \in2_data[0]~input_o  = in2_data[0];

assign \in2_data[1]~input_o  = in2_data[1];

assign \in2_data[2]~input_o  = in2_data[2];

assign \in2_data[3]~input_o  = in2_data[3];

assign \in3_data[0]~input_o  = in3_data[0];

assign \in3_data[1]~input_o  = in3_data[1];

assign \in3_data[2]~input_o  = in3_data[2];

assign \in3_data[3]~input_o  = in3_data[3];

assign \in4_data[0]~input_o  = in4_data[0];

assign \in4_data[1]~input_o  = in4_data[1];

assign \in4_data[2]~input_o  = in4_data[2];

assign \in4_data[3]~input_o  = in4_data[3];

assign \in5_data[0]~input_o  = in5_data[0];

assign \in5_data[1]~input_o  = in5_data[1];

assign \in5_data[2]~input_o  = in5_data[2];

assign \in5_data[3]~input_o  = in5_data[3];

assign \in6_data[0]~input_o  = in6_data[0];

assign \in6_data[1]~input_o  = in6_data[1];

assign \in6_data[2]~input_o  = in6_data[2];

assign \in6_data[3]~input_o  = in6_data[3];

assign \in7_data[0]~input_o  = in7_data[0];

assign \in7_data[1]~input_o  = in7_data[1];

assign \in7_data[2]~input_o  = in7_data[2];

assign \in7_data[3]~input_o  = in7_data[3];

assign \in8_data[0]~input_o  = in8_data[0];

assign \in8_data[1]~input_o  = in8_data[1];

assign \in8_data[2]~input_o  = in8_data[2];

assign \in8_data[3]~input_o  = in8_data[3];

assign \in9_data[0]~input_o  = in9_data[0];

assign \in9_data[1]~input_o  = in9_data[1];

assign \in9_data[2]~input_o  = in9_data[2];

assign \in9_data[3]~input_o  = in9_data[3];

assign \in10_data[0]~input_o  = in10_data[0];

assign \in10_data[1]~input_o  = in10_data[1];

assign \in10_data[2]~input_o  = in10_data[2];

assign \in10_data[3]~input_o  = in10_data[3];

assign \in11_data[0]~input_o  = in11_data[0];

assign \in11_data[1]~input_o  = in11_data[1];

assign \in11_data[2]~input_o  = in11_data[2];

assign \in11_data[3]~input_o  = in11_data[3];

assign \in12_data[0]~input_o  = in12_data[0];

assign \in12_data[1]~input_o  = in12_data[1];

assign \in12_data[2]~input_o  = in12_data[2];

assign \in12_data[3]~input_o  = in12_data[3];

assign \in13_data[0]~input_o  = in13_data[0];

assign \in13_data[1]~input_o  = in13_data[1];

assign \in13_data[2]~input_o  = in13_data[2];

assign \in13_data[3]~input_o  = in13_data[3];

assign \in14_data[0]~input_o  = in14_data[0];

assign \in14_data[1]~input_o  = in14_data[1];

assign \in14_data[2]~input_o  = in14_data[2];

assign \in14_data[3]~input_o  = in14_data[3];

assign \in15_data[0]~input_o  = in15_data[0];

assign \in15_data[1]~input_o  = in15_data[1];

assign \in15_data[2]~input_o  = in15_data[2];

assign \in15_data[3]~input_o  = in15_data[3];

endmodule

module CIC_CIC_cic_ii_0 (
	full_dff,
	source_valid_s,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	GND_port,
	NJQG9082,
	clk,
	in_valid,
	reset_n,
	out_ready,
	in10_data_10,
	in10_data_9,
	in10_data_8,
	in10_data_7,
	in10_data_6,
	in10_data_5,
	in10_data_4,
	in6_data_10,
	in6_data_9,
	in6_data_8,
	in6_data_7,
	in6_data_6,
	in6_data_5,
	in6_data_4,
	in14_data_10,
	in14_data_9,
	in14_data_8,
	in14_data_7,
	in14_data_6,
	in14_data_5,
	in14_data_4,
	in2_data_10,
	in2_data_9,
	in2_data_8,
	in2_data_7,
	in2_data_6,
	in2_data_5,
	in2_data_4,
	in11_data_10,
	in11_data_9,
	in11_data_8,
	in11_data_7,
	in11_data_6,
	in11_data_5,
	in11_data_4,
	in7_data_10,
	in7_data_9,
	in7_data_8,
	in7_data_7,
	in7_data_6,
	in7_data_5,
	in7_data_4,
	in15_data_10,
	in15_data_9,
	in15_data_8,
	in15_data_7,
	in15_data_6,
	in15_data_5,
	in15_data_4,
	in3_data_10,
	in3_data_9,
	in3_data_8,
	in3_data_7,
	in3_data_6,
	in3_data_5,
	in3_data_4,
	in5_data_10,
	in5_data_9,
	in5_data_8,
	in5_data_7,
	in5_data_6,
	in5_data_5,
	in5_data_4,
	in9_data_10,
	in9_data_9,
	in9_data_8,
	in9_data_7,
	in9_data_6,
	in9_data_5,
	in9_data_4,
	in13_data_10,
	in13_data_9,
	in13_data_8,
	in13_data_7,
	in13_data_6,
	in13_data_5,
	in13_data_4,
	in1_data_10,
	in1_data_9,
	in1_data_8,
	in1_data_7,
	in1_data_6,
	in1_data_5,
	in1_data_4,
	in4_data_10,
	in4_data_9,
	in4_data_8,
	in4_data_7,
	in4_data_6,
	in4_data_5,
	in4_data_4,
	in8_data_10,
	in8_data_9,
	in8_data_8,
	in8_data_7,
	in8_data_6,
	in8_data_5,
	in8_data_4,
	in12_data_10,
	in12_data_9,
	in12_data_8,
	in12_data_7,
	in12_data_6,
	in12_data_5,
	in12_data_4,
	in0_data_10,
	in0_data_9,
	in0_data_8,
	in0_data_7,
	in0_data_6,
	in0_data_5,
	in0_data_4,
	in6_data_11,
	in7_data_11,
	in5_data_11,
	in4_data_11,
	in10_data_11,
	in11_data_11,
	in9_data_11,
	in8_data_11,
	in14_data_11,
	in15_data_11,
	in13_data_11,
	in12_data_11,
	in2_data_11,
	in3_data_11,
	in1_data_11,
	in0_data_11,
	in6_data_12,
	in10_data_12,
	in14_data_12,
	in2_data_12,
	in7_data_12,
	in11_data_12,
	in15_data_12,
	in3_data_12,
	in9_data_12,
	in5_data_12,
	in13_data_12,
	in1_data_12,
	in8_data_12,
	in4_data_12,
	in12_data_12,
	in0_data_12,
	in10_data_13,
	in11_data_13,
	in9_data_13,
	in8_data_13,
	in6_data_13,
	in7_data_13,
	in5_data_13,
	in4_data_13,
	in14_data_13,
	in15_data_13,
	in13_data_13,
	in12_data_13,
	in2_data_13,
	in3_data_13,
	in1_data_13,
	in0_data_13,
	in10_data_14,
	in6_data_14,
	in14_data_14,
	in2_data_14,
	in11_data_14,
	in7_data_14,
	in15_data_14,
	in3_data_14,
	in5_data_14,
	in9_data_14,
	in13_data_14,
	in1_data_14,
	in4_data_14,
	in8_data_14,
	in12_data_14,
	in0_data_14,
	in6_data_15,
	in7_data_15,
	in5_data_15,
	in4_data_15,
	in10_data_15,
	in11_data_15,
	in9_data_15,
	in8_data_15,
	in14_data_15,
	in15_data_15,
	in13_data_15,
	in12_data_15,
	in2_data_15,
	in3_data_15,
	in1_data_15,
	in0_data_15)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	source_valid_s;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
input 	GND_port;
input 	NJQG9082;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	out_ready;
input 	in10_data_10;
input 	in10_data_9;
input 	in10_data_8;
input 	in10_data_7;
input 	in10_data_6;
input 	in10_data_5;
input 	in10_data_4;
input 	in6_data_10;
input 	in6_data_9;
input 	in6_data_8;
input 	in6_data_7;
input 	in6_data_6;
input 	in6_data_5;
input 	in6_data_4;
input 	in14_data_10;
input 	in14_data_9;
input 	in14_data_8;
input 	in14_data_7;
input 	in14_data_6;
input 	in14_data_5;
input 	in14_data_4;
input 	in2_data_10;
input 	in2_data_9;
input 	in2_data_8;
input 	in2_data_7;
input 	in2_data_6;
input 	in2_data_5;
input 	in2_data_4;
input 	in11_data_10;
input 	in11_data_9;
input 	in11_data_8;
input 	in11_data_7;
input 	in11_data_6;
input 	in11_data_5;
input 	in11_data_4;
input 	in7_data_10;
input 	in7_data_9;
input 	in7_data_8;
input 	in7_data_7;
input 	in7_data_6;
input 	in7_data_5;
input 	in7_data_4;
input 	in15_data_10;
input 	in15_data_9;
input 	in15_data_8;
input 	in15_data_7;
input 	in15_data_6;
input 	in15_data_5;
input 	in15_data_4;
input 	in3_data_10;
input 	in3_data_9;
input 	in3_data_8;
input 	in3_data_7;
input 	in3_data_6;
input 	in3_data_5;
input 	in3_data_4;
input 	in5_data_10;
input 	in5_data_9;
input 	in5_data_8;
input 	in5_data_7;
input 	in5_data_6;
input 	in5_data_5;
input 	in5_data_4;
input 	in9_data_10;
input 	in9_data_9;
input 	in9_data_8;
input 	in9_data_7;
input 	in9_data_6;
input 	in9_data_5;
input 	in9_data_4;
input 	in13_data_10;
input 	in13_data_9;
input 	in13_data_8;
input 	in13_data_7;
input 	in13_data_6;
input 	in13_data_5;
input 	in13_data_4;
input 	in1_data_10;
input 	in1_data_9;
input 	in1_data_8;
input 	in1_data_7;
input 	in1_data_6;
input 	in1_data_5;
input 	in1_data_4;
input 	in4_data_10;
input 	in4_data_9;
input 	in4_data_8;
input 	in4_data_7;
input 	in4_data_6;
input 	in4_data_5;
input 	in4_data_4;
input 	in8_data_10;
input 	in8_data_9;
input 	in8_data_8;
input 	in8_data_7;
input 	in8_data_6;
input 	in8_data_5;
input 	in8_data_4;
input 	in12_data_10;
input 	in12_data_9;
input 	in12_data_8;
input 	in12_data_7;
input 	in12_data_6;
input 	in12_data_5;
input 	in12_data_4;
input 	in0_data_10;
input 	in0_data_9;
input 	in0_data_8;
input 	in0_data_7;
input 	in0_data_6;
input 	in0_data_5;
input 	in0_data_4;
input 	in6_data_11;
input 	in7_data_11;
input 	in5_data_11;
input 	in4_data_11;
input 	in10_data_11;
input 	in11_data_11;
input 	in9_data_11;
input 	in8_data_11;
input 	in14_data_11;
input 	in15_data_11;
input 	in13_data_11;
input 	in12_data_11;
input 	in2_data_11;
input 	in3_data_11;
input 	in1_data_11;
input 	in0_data_11;
input 	in6_data_12;
input 	in10_data_12;
input 	in14_data_12;
input 	in2_data_12;
input 	in7_data_12;
input 	in11_data_12;
input 	in15_data_12;
input 	in3_data_12;
input 	in9_data_12;
input 	in5_data_12;
input 	in13_data_12;
input 	in1_data_12;
input 	in8_data_12;
input 	in4_data_12;
input 	in12_data_12;
input 	in0_data_12;
input 	in10_data_13;
input 	in11_data_13;
input 	in9_data_13;
input 	in8_data_13;
input 	in6_data_13;
input 	in7_data_13;
input 	in5_data_13;
input 	in4_data_13;
input 	in14_data_13;
input 	in15_data_13;
input 	in13_data_13;
input 	in12_data_13;
input 	in2_data_13;
input 	in3_data_13;
input 	in1_data_13;
input 	in0_data_13;
input 	in10_data_14;
input 	in6_data_14;
input 	in14_data_14;
input 	in2_data_14;
input 	in11_data_14;
input 	in7_data_14;
input 	in15_data_14;
input 	in3_data_14;
input 	in5_data_14;
input 	in9_data_14;
input 	in13_data_14;
input 	in1_data_14;
input 	in4_data_14;
input 	in8_data_14;
input 	in12_data_14;
input 	in0_data_14;
input 	in6_data_15;
input 	in7_data_15;
input 	in5_data_15;
input 	in4_data_15;
input 	in10_data_15;
input 	in11_data_15;
input 	in9_data_15;
input 	in8_data_15;
input 	in14_data_15;
input 	in15_data_15;
input 	in13_data_15;
input 	in12_data_15;
input 	in2_data_15;
input 	in3_data_15;
input 	in1_data_15;
input 	in0_data_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;


CIC_alt_cic_core core(
	.full_dff(full_dff),
	.q_b_0(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_8(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_9(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_10(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_11(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_12(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_13(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_14(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_15(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.source_valid_s(source_valid_s),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.GND_port(GND_port),
	.clk(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.out_ready(out_ready),
	.in10_data_10(in10_data_10),
	.in10_data_9(in10_data_9),
	.in10_data_8(in10_data_8),
	.in10_data_7(in10_data_7),
	.in10_data_6(in10_data_6),
	.in10_data_5(in10_data_5),
	.in10_data_4(in10_data_4),
	.in6_data_10(in6_data_10),
	.in6_data_9(in6_data_9),
	.in6_data_8(in6_data_8),
	.in6_data_7(in6_data_7),
	.in6_data_6(in6_data_6),
	.in6_data_5(in6_data_5),
	.in6_data_4(in6_data_4),
	.in14_data_10(in14_data_10),
	.in14_data_9(in14_data_9),
	.in14_data_8(in14_data_8),
	.in14_data_7(in14_data_7),
	.in14_data_6(in14_data_6),
	.in14_data_5(in14_data_5),
	.in14_data_4(in14_data_4),
	.in2_data_10(in2_data_10),
	.in2_data_9(in2_data_9),
	.in2_data_8(in2_data_8),
	.in2_data_7(in2_data_7),
	.in2_data_6(in2_data_6),
	.in2_data_5(in2_data_5),
	.in2_data_4(in2_data_4),
	.in11_data_10(in11_data_10),
	.in11_data_9(in11_data_9),
	.in11_data_8(in11_data_8),
	.in11_data_7(in11_data_7),
	.in11_data_6(in11_data_6),
	.in11_data_5(in11_data_5),
	.in11_data_4(in11_data_4),
	.in7_data_10(in7_data_10),
	.in7_data_9(in7_data_9),
	.in7_data_8(in7_data_8),
	.in7_data_7(in7_data_7),
	.in7_data_6(in7_data_6),
	.in7_data_5(in7_data_5),
	.in7_data_4(in7_data_4),
	.in15_data_10(in15_data_10),
	.in15_data_9(in15_data_9),
	.in15_data_8(in15_data_8),
	.in15_data_7(in15_data_7),
	.in15_data_6(in15_data_6),
	.in15_data_5(in15_data_5),
	.in15_data_4(in15_data_4),
	.in3_data_10(in3_data_10),
	.in3_data_9(in3_data_9),
	.in3_data_8(in3_data_8),
	.in3_data_7(in3_data_7),
	.in3_data_6(in3_data_6),
	.in3_data_5(in3_data_5),
	.in3_data_4(in3_data_4),
	.in5_data_10(in5_data_10),
	.in5_data_9(in5_data_9),
	.in5_data_8(in5_data_8),
	.in5_data_7(in5_data_7),
	.in5_data_6(in5_data_6),
	.in5_data_5(in5_data_5),
	.in5_data_4(in5_data_4),
	.in9_data_10(in9_data_10),
	.in9_data_9(in9_data_9),
	.in9_data_8(in9_data_8),
	.in9_data_7(in9_data_7),
	.in9_data_6(in9_data_6),
	.in9_data_5(in9_data_5),
	.in9_data_4(in9_data_4),
	.in13_data_10(in13_data_10),
	.in13_data_9(in13_data_9),
	.in13_data_8(in13_data_8),
	.in13_data_7(in13_data_7),
	.in13_data_6(in13_data_6),
	.in13_data_5(in13_data_5),
	.in13_data_4(in13_data_4),
	.in1_data_10(in1_data_10),
	.in1_data_9(in1_data_9),
	.in1_data_8(in1_data_8),
	.in1_data_7(in1_data_7),
	.in1_data_6(in1_data_6),
	.in1_data_5(in1_data_5),
	.in1_data_4(in1_data_4),
	.in4_data_10(in4_data_10),
	.in4_data_9(in4_data_9),
	.in4_data_8(in4_data_8),
	.in4_data_7(in4_data_7),
	.in4_data_6(in4_data_6),
	.in4_data_5(in4_data_5),
	.in4_data_4(in4_data_4),
	.in8_data_10(in8_data_10),
	.in8_data_9(in8_data_9),
	.in8_data_8(in8_data_8),
	.in8_data_7(in8_data_7),
	.in8_data_6(in8_data_6),
	.in8_data_5(in8_data_5),
	.in8_data_4(in8_data_4),
	.in12_data_10(in12_data_10),
	.in12_data_9(in12_data_9),
	.in12_data_8(in12_data_8),
	.in12_data_7(in12_data_7),
	.in12_data_6(in12_data_6),
	.in12_data_5(in12_data_5),
	.in12_data_4(in12_data_4),
	.in0_data_10(in0_data_10),
	.in0_data_9(in0_data_9),
	.in0_data_8(in0_data_8),
	.in0_data_7(in0_data_7),
	.in0_data_6(in0_data_6),
	.in0_data_5(in0_data_5),
	.in0_data_4(in0_data_4),
	.in6_data_11(in6_data_11),
	.in7_data_11(in7_data_11),
	.in5_data_11(in5_data_11),
	.in4_data_11(in4_data_11),
	.in10_data_11(in10_data_11),
	.in11_data_11(in11_data_11),
	.in9_data_11(in9_data_11),
	.in8_data_11(in8_data_11),
	.in14_data_11(in14_data_11),
	.in15_data_11(in15_data_11),
	.in13_data_11(in13_data_11),
	.in12_data_11(in12_data_11),
	.in2_data_11(in2_data_11),
	.in3_data_11(in3_data_11),
	.in1_data_11(in1_data_11),
	.in0_data_11(in0_data_11),
	.in6_data_12(in6_data_12),
	.in10_data_12(in10_data_12),
	.in14_data_12(in14_data_12),
	.in2_data_12(in2_data_12),
	.in7_data_12(in7_data_12),
	.in11_data_12(in11_data_12),
	.in15_data_12(in15_data_12),
	.in3_data_12(in3_data_12),
	.in9_data_12(in9_data_12),
	.in5_data_12(in5_data_12),
	.in13_data_12(in13_data_12),
	.in1_data_12(in1_data_12),
	.in8_data_12(in8_data_12),
	.in4_data_12(in4_data_12),
	.in12_data_12(in12_data_12),
	.in0_data_12(in0_data_12),
	.in10_data_13(in10_data_13),
	.in11_data_13(in11_data_13),
	.in9_data_13(in9_data_13),
	.in8_data_13(in8_data_13),
	.in6_data_13(in6_data_13),
	.in7_data_13(in7_data_13),
	.in5_data_13(in5_data_13),
	.in4_data_13(in4_data_13),
	.in14_data_13(in14_data_13),
	.in15_data_13(in15_data_13),
	.in13_data_13(in13_data_13),
	.in12_data_13(in12_data_13),
	.in2_data_13(in2_data_13),
	.in3_data_13(in3_data_13),
	.in1_data_13(in1_data_13),
	.in0_data_13(in0_data_13),
	.in10_data_14(in10_data_14),
	.in6_data_14(in6_data_14),
	.in14_data_14(in14_data_14),
	.in2_data_14(in2_data_14),
	.in11_data_14(in11_data_14),
	.in7_data_14(in7_data_14),
	.in15_data_14(in15_data_14),
	.in3_data_14(in3_data_14),
	.in5_data_14(in5_data_14),
	.in9_data_14(in9_data_14),
	.in13_data_14(in13_data_14),
	.in1_data_14(in1_data_14),
	.in4_data_14(in4_data_14),
	.in8_data_14(in8_data_14),
	.in12_data_14(in12_data_14),
	.in0_data_14(in0_data_14),
	.in6_data_15(in6_data_15),
	.in7_data_15(in7_data_15),
	.in5_data_15(in5_data_15),
	.in4_data_15(in4_data_15),
	.in10_data_15(in10_data_15),
	.in11_data_15(in11_data_15),
	.in9_data_15(in9_data_15),
	.in8_data_15(in8_data_15),
	.in14_data_15(in14_data_15),
	.in15_data_15(in15_data_15),
	.in13_data_15(in13_data_15),
	.in12_data_15(in12_data_15),
	.in2_data_15(in2_data_15),
	.in3_data_15(in3_data_15),
	.in1_data_15(in1_data_15),
	.in0_data_15(in0_data_15));

cycloneive_lcell_comb \out_data[0] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_0),
	.cout());
defparam \out_data[0] .lut_mask = 16'hAAFF;
defparam \out_data[0] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[1] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_1),
	.cout());
defparam \out_data[1] .lut_mask = 16'hAAFF;
defparam \out_data[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[2] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_2),
	.cout());
defparam \out_data[2] .lut_mask = 16'hAAFF;
defparam \out_data[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[3] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_3),
	.cout());
defparam \out_data[3] .lut_mask = 16'hAAFF;
defparam \out_data[3] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[4] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_4),
	.cout());
defparam \out_data[4] .lut_mask = 16'hAAFF;
defparam \out_data[4] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[5] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5] .lut_mask = 16'hAAFF;
defparam \out_data[5] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[6] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_6),
	.cout());
defparam \out_data[6] .lut_mask = 16'hAAFF;
defparam \out_data[6] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[7] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_7),
	.cout());
defparam \out_data[7] .lut_mask = 16'hAAFF;
defparam \out_data[7] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[8] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_8),
	.cout());
defparam \out_data[8] .lut_mask = 16'hAAFF;
defparam \out_data[8] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[9] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_9),
	.cout());
defparam \out_data[9] .lut_mask = 16'hAAFF;
defparam \out_data[9] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[10] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_10),
	.cout());
defparam \out_data[10] .lut_mask = 16'hAAFF;
defparam \out_data[10] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[11] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_11),
	.cout());
defparam \out_data[11] .lut_mask = 16'hAAFF;
defparam \out_data[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[12] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_12),
	.cout());
defparam \out_data[12] .lut_mask = 16'hAAFF;
defparam \out_data[12] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[13] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_13),
	.cout());
defparam \out_data[13] .lut_mask = 16'hAAFF;
defparam \out_data[13] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[14] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_14),
	.cout());
defparam \out_data[14] .lut_mask = 16'hAAFF;
defparam \out_data[14] .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_data[15] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_15),
	.cout());
defparam \out_data[15] .lut_mask = 16'hAAFF;
defparam \out_data[15] .sum_lutc_input = "datac";

endmodule

module CIC_alt_cic_core (
	full_dff,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	source_valid_s,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	GND_port,
	clk,
	in_valid,
	reset_n,
	out_ready,
	in10_data_10,
	in10_data_9,
	in10_data_8,
	in10_data_7,
	in10_data_6,
	in10_data_5,
	in10_data_4,
	in6_data_10,
	in6_data_9,
	in6_data_8,
	in6_data_7,
	in6_data_6,
	in6_data_5,
	in6_data_4,
	in14_data_10,
	in14_data_9,
	in14_data_8,
	in14_data_7,
	in14_data_6,
	in14_data_5,
	in14_data_4,
	in2_data_10,
	in2_data_9,
	in2_data_8,
	in2_data_7,
	in2_data_6,
	in2_data_5,
	in2_data_4,
	in11_data_10,
	in11_data_9,
	in11_data_8,
	in11_data_7,
	in11_data_6,
	in11_data_5,
	in11_data_4,
	in7_data_10,
	in7_data_9,
	in7_data_8,
	in7_data_7,
	in7_data_6,
	in7_data_5,
	in7_data_4,
	in15_data_10,
	in15_data_9,
	in15_data_8,
	in15_data_7,
	in15_data_6,
	in15_data_5,
	in15_data_4,
	in3_data_10,
	in3_data_9,
	in3_data_8,
	in3_data_7,
	in3_data_6,
	in3_data_5,
	in3_data_4,
	in5_data_10,
	in5_data_9,
	in5_data_8,
	in5_data_7,
	in5_data_6,
	in5_data_5,
	in5_data_4,
	in9_data_10,
	in9_data_9,
	in9_data_8,
	in9_data_7,
	in9_data_6,
	in9_data_5,
	in9_data_4,
	in13_data_10,
	in13_data_9,
	in13_data_8,
	in13_data_7,
	in13_data_6,
	in13_data_5,
	in13_data_4,
	in1_data_10,
	in1_data_9,
	in1_data_8,
	in1_data_7,
	in1_data_6,
	in1_data_5,
	in1_data_4,
	in4_data_10,
	in4_data_9,
	in4_data_8,
	in4_data_7,
	in4_data_6,
	in4_data_5,
	in4_data_4,
	in8_data_10,
	in8_data_9,
	in8_data_8,
	in8_data_7,
	in8_data_6,
	in8_data_5,
	in8_data_4,
	in12_data_10,
	in12_data_9,
	in12_data_8,
	in12_data_7,
	in12_data_6,
	in12_data_5,
	in12_data_4,
	in0_data_10,
	in0_data_9,
	in0_data_8,
	in0_data_7,
	in0_data_6,
	in0_data_5,
	in0_data_4,
	in6_data_11,
	in7_data_11,
	in5_data_11,
	in4_data_11,
	in10_data_11,
	in11_data_11,
	in9_data_11,
	in8_data_11,
	in14_data_11,
	in15_data_11,
	in13_data_11,
	in12_data_11,
	in2_data_11,
	in3_data_11,
	in1_data_11,
	in0_data_11,
	in6_data_12,
	in10_data_12,
	in14_data_12,
	in2_data_12,
	in7_data_12,
	in11_data_12,
	in15_data_12,
	in3_data_12,
	in9_data_12,
	in5_data_12,
	in13_data_12,
	in1_data_12,
	in8_data_12,
	in4_data_12,
	in12_data_12,
	in0_data_12,
	in10_data_13,
	in11_data_13,
	in9_data_13,
	in8_data_13,
	in6_data_13,
	in7_data_13,
	in5_data_13,
	in4_data_13,
	in14_data_13,
	in15_data_13,
	in13_data_13,
	in12_data_13,
	in2_data_13,
	in3_data_13,
	in1_data_13,
	in0_data_13,
	in10_data_14,
	in6_data_14,
	in14_data_14,
	in2_data_14,
	in11_data_14,
	in7_data_14,
	in15_data_14,
	in3_data_14,
	in5_data_14,
	in9_data_14,
	in13_data_14,
	in1_data_14,
	in4_data_14,
	in8_data_14,
	in12_data_14,
	in0_data_14,
	in6_data_15,
	in7_data_15,
	in5_data_15,
	in4_data_15,
	in10_data_15,
	in11_data_15,
	in9_data_15,
	in8_data_15,
	in14_data_15,
	in15_data_15,
	in13_data_15,
	in12_data_15,
	in2_data_15,
	in3_data_15,
	in1_data_15,
	in0_data_15)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	source_valid_s;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
input 	GND_port;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	out_ready;
input 	in10_data_10;
input 	in10_data_9;
input 	in10_data_8;
input 	in10_data_7;
input 	in10_data_6;
input 	in10_data_5;
input 	in10_data_4;
input 	in6_data_10;
input 	in6_data_9;
input 	in6_data_8;
input 	in6_data_7;
input 	in6_data_6;
input 	in6_data_5;
input 	in6_data_4;
input 	in14_data_10;
input 	in14_data_9;
input 	in14_data_8;
input 	in14_data_7;
input 	in14_data_6;
input 	in14_data_5;
input 	in14_data_4;
input 	in2_data_10;
input 	in2_data_9;
input 	in2_data_8;
input 	in2_data_7;
input 	in2_data_6;
input 	in2_data_5;
input 	in2_data_4;
input 	in11_data_10;
input 	in11_data_9;
input 	in11_data_8;
input 	in11_data_7;
input 	in11_data_6;
input 	in11_data_5;
input 	in11_data_4;
input 	in7_data_10;
input 	in7_data_9;
input 	in7_data_8;
input 	in7_data_7;
input 	in7_data_6;
input 	in7_data_5;
input 	in7_data_4;
input 	in15_data_10;
input 	in15_data_9;
input 	in15_data_8;
input 	in15_data_7;
input 	in15_data_6;
input 	in15_data_5;
input 	in15_data_4;
input 	in3_data_10;
input 	in3_data_9;
input 	in3_data_8;
input 	in3_data_7;
input 	in3_data_6;
input 	in3_data_5;
input 	in3_data_4;
input 	in5_data_10;
input 	in5_data_9;
input 	in5_data_8;
input 	in5_data_7;
input 	in5_data_6;
input 	in5_data_5;
input 	in5_data_4;
input 	in9_data_10;
input 	in9_data_9;
input 	in9_data_8;
input 	in9_data_7;
input 	in9_data_6;
input 	in9_data_5;
input 	in9_data_4;
input 	in13_data_10;
input 	in13_data_9;
input 	in13_data_8;
input 	in13_data_7;
input 	in13_data_6;
input 	in13_data_5;
input 	in13_data_4;
input 	in1_data_10;
input 	in1_data_9;
input 	in1_data_8;
input 	in1_data_7;
input 	in1_data_6;
input 	in1_data_5;
input 	in1_data_4;
input 	in4_data_10;
input 	in4_data_9;
input 	in4_data_8;
input 	in4_data_7;
input 	in4_data_6;
input 	in4_data_5;
input 	in4_data_4;
input 	in8_data_10;
input 	in8_data_9;
input 	in8_data_8;
input 	in8_data_7;
input 	in8_data_6;
input 	in8_data_5;
input 	in8_data_4;
input 	in12_data_10;
input 	in12_data_9;
input 	in12_data_8;
input 	in12_data_7;
input 	in12_data_6;
input 	in12_data_5;
input 	in12_data_4;
input 	in0_data_10;
input 	in0_data_9;
input 	in0_data_8;
input 	in0_data_7;
input 	in0_data_6;
input 	in0_data_5;
input 	in0_data_4;
input 	in6_data_11;
input 	in7_data_11;
input 	in5_data_11;
input 	in4_data_11;
input 	in10_data_11;
input 	in11_data_11;
input 	in9_data_11;
input 	in8_data_11;
input 	in14_data_11;
input 	in15_data_11;
input 	in13_data_11;
input 	in12_data_11;
input 	in2_data_11;
input 	in3_data_11;
input 	in1_data_11;
input 	in0_data_11;
input 	in6_data_12;
input 	in10_data_12;
input 	in14_data_12;
input 	in2_data_12;
input 	in7_data_12;
input 	in11_data_12;
input 	in15_data_12;
input 	in3_data_12;
input 	in9_data_12;
input 	in5_data_12;
input 	in13_data_12;
input 	in1_data_12;
input 	in8_data_12;
input 	in4_data_12;
input 	in12_data_12;
input 	in0_data_12;
input 	in10_data_13;
input 	in11_data_13;
input 	in9_data_13;
input 	in8_data_13;
input 	in6_data_13;
input 	in7_data_13;
input 	in5_data_13;
input 	in4_data_13;
input 	in14_data_13;
input 	in15_data_13;
input 	in13_data_13;
input 	in12_data_13;
input 	in2_data_13;
input 	in3_data_13;
input 	in1_data_13;
input 	in0_data_13;
input 	in10_data_14;
input 	in6_data_14;
input 	in14_data_14;
input 	in2_data_14;
input 	in11_data_14;
input 	in7_data_14;
input 	in15_data_14;
input 	in3_data_14;
input 	in5_data_14;
input 	in9_data_14;
input 	in13_data_14;
input 	in1_data_14;
input 	in4_data_14;
input 	in8_data_14;
input 	in12_data_14;
input 	in0_data_14;
input 	in6_data_15;
input 	in7_data_15;
input 	in5_data_15;
input 	in4_data_15;
input 	in10_data_15;
input 	in11_data_15;
input 	in9_data_15;
input 	in8_data_15;
input 	in14_data_15;
input 	in15_data_15;
input 	in13_data_15;
input 	in12_data_15;
input 	in2_data_15;
input 	in3_data_15;
input 	in1_data_15;
input 	in0_data_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \input_sink|sink_FIFO|auto_generated|dffe_nae~q ;
wire \output_source_1|source_FIFO|auto_generated|dffe_af~q ;
wire \dec_mul|state[0]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[1]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[2]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[3]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[4]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[5]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[6]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[7]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[8]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[9]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[10]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[11]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[12]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[13]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[14]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[15]~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout[16]~q ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[170] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[169] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[168] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[167] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[166] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[165] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[164] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[106] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[105] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[104] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[103] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[102] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[101] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[100] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[234] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[233] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[232] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[231] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[230] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[229] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[228] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[42] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[41] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[40] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[39] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[38] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[37] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[36] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[186] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[185] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[184] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[183] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[182] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[181] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[180] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[122] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[121] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[120] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[119] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[118] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[117] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[116] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[250] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[249] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[248] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[247] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[246] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[245] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[244] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[58] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[57] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[56] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[55] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[54] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[53] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[52] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[90] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[89] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[88] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[87] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[86] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[85] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[84] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[154] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[153] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[152] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[151] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[150] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[149] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[148] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[218] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[217] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[216] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[215] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[214] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[213] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[212] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[74] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[73] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[72] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[71] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[70] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[69] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[68] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[138] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[137] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[136] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[135] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[134] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[133] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[132] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[202] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[201] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[200] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[199] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[198] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[197] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[196] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[107] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[123] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[91] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[75] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[171] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[187] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[155] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[139] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[235] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[251] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[219] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[203] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[43] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[59] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[108] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[172] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[236] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[44] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[124] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[188] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[252] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[60] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[156] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[92] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[220] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[140] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[76] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[204] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[173] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[189] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[157] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[141] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[109] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[125] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[93] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[77] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[237] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[253] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[221] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[205] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[45] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[61] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[174] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[110] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[238] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[46] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[190] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[126] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[254] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[62] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[94] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[158] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[222] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[78] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[142] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[206] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[111] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[127] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[95] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[79] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[175] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[191] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[159] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[143] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[239] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[255] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[223] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[207] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[47] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[63] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \avalon_controller|sink_ready_ctrl~2_combout ;
wire \avalon_controller|stall_reg~q ;
wire \dec_mul|stage_diff[0].auk_dsp_diff|dout_valid~q ;
wire \dec_mul|channel_out_int[0]~q ;
wire \dec_mul|channel_out_int[1]~q ;
wire \dec_mul|channel_out_int[2]~q ;
wire \dec_mul|channel_out_int[3]~q ;
wire \avalon_controller|ready_FIFO|usedw_process~0_combout ;


CIC_alt_cic_dec_miso dec_mul(
	.state_0(\dec_mul|state[0]~q ),
	.dout_1(\dec_mul|stage_diff[0].auk_dsp_diff|dout[1]~q ),
	.dout_2(\dec_mul|stage_diff[0].auk_dsp_diff|dout[2]~q ),
	.dout_3(\dec_mul|stage_diff[0].auk_dsp_diff|dout[3]~q ),
	.dout_4(\dec_mul|stage_diff[0].auk_dsp_diff|dout[4]~q ),
	.dout_5(\dec_mul|stage_diff[0].auk_dsp_diff|dout[5]~q ),
	.dout_6(\dec_mul|stage_diff[0].auk_dsp_diff|dout[6]~q ),
	.dout_7(\dec_mul|stage_diff[0].auk_dsp_diff|dout[7]~q ),
	.dout_8(\dec_mul|stage_diff[0].auk_dsp_diff|dout[8]~q ),
	.dout_9(\dec_mul|stage_diff[0].auk_dsp_diff|dout[9]~q ),
	.dout_10(\dec_mul|stage_diff[0].auk_dsp_diff|dout[10]~q ),
	.dout_11(\dec_mul|stage_diff[0].auk_dsp_diff|dout[11]~q ),
	.dout_12(\dec_mul|stage_diff[0].auk_dsp_diff|dout[12]~q ),
	.dout_13(\dec_mul|stage_diff[0].auk_dsp_diff|dout[13]~q ),
	.dout_14(\dec_mul|stage_diff[0].auk_dsp_diff|dout[14]~q ),
	.dout_15(\dec_mul|stage_diff[0].auk_dsp_diff|dout[15]~q ),
	.dout_16(\dec_mul|stage_diff[0].auk_dsp_diff|dout[16]~q ),
	.q_b_170(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[170] ),
	.q_b_169(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[169] ),
	.q_b_168(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[168] ),
	.q_b_167(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[167] ),
	.q_b_166(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[166] ),
	.q_b_165(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[165] ),
	.q_b_164(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[164] ),
	.q_b_106(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[106] ),
	.q_b_105(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[105] ),
	.q_b_104(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[104] ),
	.q_b_103(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[103] ),
	.q_b_102(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[102] ),
	.q_b_101(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[101] ),
	.q_b_100(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[100] ),
	.q_b_234(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[234] ),
	.q_b_233(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[233] ),
	.q_b_232(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[232] ),
	.q_b_231(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[231] ),
	.q_b_230(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[230] ),
	.q_b_229(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[229] ),
	.q_b_228(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[228] ),
	.q_b_42(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[42] ),
	.q_b_41(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[41] ),
	.q_b_40(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[40] ),
	.q_b_39(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[39] ),
	.q_b_38(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[38] ),
	.q_b_37(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[37] ),
	.q_b_36(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[36] ),
	.q_b_186(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[186] ),
	.q_b_185(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[185] ),
	.q_b_184(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[184] ),
	.q_b_183(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[183] ),
	.q_b_182(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[182] ),
	.q_b_181(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[181] ),
	.q_b_180(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[180] ),
	.q_b_122(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[122] ),
	.q_b_121(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[121] ),
	.q_b_120(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[120] ),
	.q_b_119(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[119] ),
	.q_b_118(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[118] ),
	.q_b_117(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[117] ),
	.q_b_116(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[116] ),
	.q_b_250(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[250] ),
	.q_b_249(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[249] ),
	.q_b_248(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[248] ),
	.q_b_247(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[247] ),
	.q_b_246(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[246] ),
	.q_b_245(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[245] ),
	.q_b_244(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[244] ),
	.q_b_58(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[58] ),
	.q_b_57(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[57] ),
	.q_b_56(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[56] ),
	.q_b_55(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[55] ),
	.q_b_54(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[54] ),
	.q_b_53(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[53] ),
	.q_b_52(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[52] ),
	.q_b_90(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[90] ),
	.q_b_89(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[89] ),
	.q_b_88(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[88] ),
	.q_b_87(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[87] ),
	.q_b_86(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[86] ),
	.q_b_85(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[85] ),
	.q_b_84(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[84] ),
	.q_b_154(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[154] ),
	.q_b_153(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[153] ),
	.q_b_152(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[152] ),
	.q_b_151(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[151] ),
	.q_b_150(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[150] ),
	.q_b_149(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[149] ),
	.q_b_148(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[148] ),
	.q_b_218(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[218] ),
	.q_b_217(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[217] ),
	.q_b_216(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[216] ),
	.q_b_215(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[215] ),
	.q_b_214(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[214] ),
	.q_b_213(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[213] ),
	.q_b_212(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[212] ),
	.q_b_26(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_25(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_24(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_23(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_22(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_21(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_20(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_74(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[74] ),
	.q_b_73(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[73] ),
	.q_b_72(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[72] ),
	.q_b_71(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[71] ),
	.q_b_70(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[70] ),
	.q_b_69(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[69] ),
	.q_b_68(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[68] ),
	.q_b_138(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[138] ),
	.q_b_137(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[137] ),
	.q_b_136(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[136] ),
	.q_b_135(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[135] ),
	.q_b_134(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[134] ),
	.q_b_133(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[133] ),
	.q_b_132(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[132] ),
	.q_b_202(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[202] ),
	.q_b_201(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[201] ),
	.q_b_200(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[200] ),
	.q_b_199(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[199] ),
	.q_b_198(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[198] ),
	.q_b_197(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[197] ),
	.q_b_196(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[196] ),
	.q_b_10(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_9(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_8(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_7(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_6(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_5(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_4(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_107(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[107] ),
	.q_b_123(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[123] ),
	.q_b_91(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[91] ),
	.q_b_75(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[75] ),
	.q_b_171(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[171] ),
	.q_b_187(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[187] ),
	.q_b_155(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[155] ),
	.q_b_139(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[139] ),
	.q_b_235(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[235] ),
	.q_b_251(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[251] ),
	.q_b_219(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[219] ),
	.q_b_203(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[203] ),
	.q_b_43(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[43] ),
	.q_b_59(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[59] ),
	.q_b_27(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_11(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_108(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[108] ),
	.q_b_172(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[172] ),
	.q_b_236(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[236] ),
	.q_b_44(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[44] ),
	.q_b_124(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[124] ),
	.q_b_188(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[188] ),
	.q_b_252(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[252] ),
	.q_b_60(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[60] ),
	.q_b_156(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[156] ),
	.q_b_92(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[92] ),
	.q_b_220(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[220] ),
	.q_b_28(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_140(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[140] ),
	.q_b_76(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[76] ),
	.q_b_204(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[204] ),
	.q_b_12(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_173(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[173] ),
	.q_b_189(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[189] ),
	.q_b_157(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[157] ),
	.q_b_141(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[141] ),
	.q_b_109(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[109] ),
	.q_b_125(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[125] ),
	.q_b_93(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[93] ),
	.q_b_77(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[77] ),
	.q_b_237(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[237] ),
	.q_b_253(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[253] ),
	.q_b_221(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[221] ),
	.q_b_205(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[205] ),
	.q_b_45(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[45] ),
	.q_b_61(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[61] ),
	.q_b_29(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_13(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_174(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[174] ),
	.q_b_110(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[110] ),
	.q_b_238(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[238] ),
	.q_b_46(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[46] ),
	.q_b_190(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[190] ),
	.q_b_126(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[126] ),
	.q_b_254(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[254] ),
	.q_b_62(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[62] ),
	.q_b_94(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[94] ),
	.q_b_158(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[158] ),
	.q_b_222(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[222] ),
	.q_b_30(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_78(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[78] ),
	.q_b_142(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[142] ),
	.q_b_206(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[206] ),
	.q_b_14(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_111(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[111] ),
	.q_b_127(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[127] ),
	.q_b_95(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[95] ),
	.q_b_79(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[79] ),
	.q_b_175(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[175] ),
	.q_b_191(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[191] ),
	.q_b_159(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[159] ),
	.q_b_143(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[143] ),
	.q_b_239(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[239] ),
	.q_b_255(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[255] ),
	.q_b_223(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[223] ),
	.q_b_207(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[207] ),
	.q_b_47(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[47] ),
	.q_b_63(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[63] ),
	.q_b_31(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.q_b_15(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.stall_reg(\avalon_controller|stall_reg~q ),
	.dout_valid(\dec_mul|stage_diff[0].auk_dsp_diff|dout_valid~q ),
	.channel_out_int_0(\dec_mul|channel_out_int[0]~q ),
	.channel_out_int_1(\dec_mul|channel_out_int[1]~q ),
	.channel_out_int_2(\dec_mul|channel_out_int[2]~q ),
	.channel_out_int_3(\dec_mul|channel_out_int[3]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_avalon_streaming_controller avalon_controller(
	.dffe_nae(\input_sink|sink_FIFO|auto_generated|dffe_nae~q ),
	.dffe_af(\output_source_1|source_FIFO|auto_generated|dffe_af~q ),
	.sink_ready_ctrl(\avalon_controller|sink_ready_ctrl~2_combout ),
	.stall_reg1(\avalon_controller|stall_reg~q ),
	.usedw_process(\avalon_controller|ready_FIFO|usedw_process~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_avalon_streaming_source output_source_1(
	.at_source_data({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.source_valid_s1(source_valid_s),
	.at_source_channel({q_b_19,q_b_18,q_b_17,q_b_16}),
	.dffe_af(\output_source_1|source_FIFO|auto_generated|dffe_af~q ),
	.state_0(\dec_mul|state[0]~q ),
	.data({\dec_mul|stage_diff[0].auk_dsp_diff|dout[16]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[15]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[14]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[13]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[12]~q ,
\dec_mul|stage_diff[0].auk_dsp_diff|dout[11]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[10]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[9]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[8]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[7]~q ,
\dec_mul|stage_diff[0].auk_dsp_diff|dout[6]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[5]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[4]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[3]~q ,\dec_mul|stage_diff[0].auk_dsp_diff|dout[2]~q ,
\dec_mul|stage_diff[0].auk_dsp_diff|dout[1]~q }),
	.stall_reg(\avalon_controller|stall_reg~q ),
	.dout_valid(\dec_mul|stage_diff[0].auk_dsp_diff|dout_valid~q ),
	.data_count({\dec_mul|channel_out_int[3]~q ,\dec_mul|channel_out_int[2]~q ,\dec_mul|channel_out_int[1]~q ,\dec_mul|channel_out_int[0]~q }),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n),
	.out_ready(out_ready));

CIC_auk_dspip_avalon_streaming_sink input_sink(
	.full_dff(full_dff),
	.dffe_nae(\input_sink|sink_FIFO|auto_generated|dffe_nae~q ),
	.dffe_af(\output_source_1|source_FIFO|auto_generated|dffe_af~q ),
	.data({\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[255] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[254] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[253] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[252] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[251] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[250] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[249] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[248] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[247] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[246] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[245] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[244] ,
data_unconnected_wire_243,data_unconnected_wire_242,data_unconnected_wire_241,data_unconnected_wire_240,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[239] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[238] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[237] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[236] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[235] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[234] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[233] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[232] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[231] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[230] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[229] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[228] ,data_unconnected_wire_227,data_unconnected_wire_226,data_unconnected_wire_225,data_unconnected_wire_224,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[223] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[222] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[221] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[220] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[219] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[218] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[217] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[216] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[215] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[214] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[213] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[212] ,
data_unconnected_wire_211,data_unconnected_wire_210,data_unconnected_wire_209,data_unconnected_wire_208,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[207] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[206] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[205] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[204] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[203] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[202] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[201] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[200] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[199] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[198] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[197] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[196] ,data_unconnected_wire_195,data_unconnected_wire_194,data_unconnected_wire_193,data_unconnected_wire_192,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[191] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[190] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[189] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[188] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[187] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[186] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[185] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[184] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[183] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[182] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[181] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[180] ,
data_unconnected_wire_179,data_unconnected_wire_178,data_unconnected_wire_177,data_unconnected_wire_176,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[175] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[174] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[173] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[172] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[171] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[170] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[169] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[168] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[167] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[166] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[165] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[164] ,data_unconnected_wire_163,data_unconnected_wire_162,data_unconnected_wire_161,data_unconnected_wire_160,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[159] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[158] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[157] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[156] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[155] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[154] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[153] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[152] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[151] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[150] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[149] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[148] ,
data_unconnected_wire_147,data_unconnected_wire_146,data_unconnected_wire_145,data_unconnected_wire_144,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[143] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[142] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[141] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[140] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[139] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[138] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[137] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[136] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[135] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[134] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[133] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[132] ,data_unconnected_wire_131,data_unconnected_wire_130,data_unconnected_wire_129,data_unconnected_wire_128,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[127] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[126] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[125] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[124] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[123] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[122] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[121] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[120] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[119] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[118] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[117] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[116] ,
data_unconnected_wire_115,data_unconnected_wire_114,data_unconnected_wire_113,data_unconnected_wire_112,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[111] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[110] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[109] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[108] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[107] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[106] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[105] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[104] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[103] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[102] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[101] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[100] ,data_unconnected_wire_99,data_unconnected_wire_98,data_unconnected_wire_97,data_unconnected_wire_96,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[95] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[94] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[93] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[92] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[91] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[90] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[89] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[88] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[87] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[86] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[85] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[84] ,
data_unconnected_wire_83,data_unconnected_wire_82,data_unconnected_wire_81,data_unconnected_wire_80,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[79] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[78] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[77] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[76] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[75] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[74] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[73] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[72] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[71] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[70] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[69] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[68] ,data_unconnected_wire_67,data_unconnected_wire_66,data_unconnected_wire_65,data_unconnected_wire_64,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[63] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[62] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[61] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[60] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[59] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[58] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[57] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[56] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[55] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[54] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[53] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[52] ,
data_unconnected_wire_51,data_unconnected_wire_50,data_unconnected_wire_49,data_unconnected_wire_48,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[47] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[46] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[45] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[44] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[43] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[42] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[41] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[40] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[39] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[38] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[37] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[36] ,data_unconnected_wire_35,data_unconnected_wire_34,data_unconnected_wire_33,data_unconnected_wire_32,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[31] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[30] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[29] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[28] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[27] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[26] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[25] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[24] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[23] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,
data_unconnected_wire_19,data_unconnected_wire_18,data_unconnected_wire_17,data_unconnected_wire_16,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,data_unconnected_wire_3,data_unconnected_wire_2,data_unconnected_wire_1,data_unconnected_wire_0}),
	.sink_ready_ctrl(\avalon_controller|sink_ready_ctrl~2_combout ),
	.usedw_process(\avalon_controller|ready_FIFO|usedw_process~0_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.at_sink_data({in15_data_15,in15_data_14,in15_data_13,in15_data_12,in15_data_11,in15_data_10,in15_data_9,in15_data_8,in15_data_7,in15_data_6,in15_data_5,in15_data_4,gnd,gnd,gnd,gnd,in14_data_15,in14_data_14,in14_data_13,in14_data_12,in14_data_11,in14_data_10,in14_data_9,in14_data_8,in14_data_7,
in14_data_6,in14_data_5,in14_data_4,gnd,gnd,gnd,gnd,in13_data_15,in13_data_14,in13_data_13,in13_data_12,in13_data_11,in13_data_10,in13_data_9,in13_data_8,in13_data_7,in13_data_6,in13_data_5,in13_data_4,gnd,gnd,gnd,gnd,in12_data_15,in12_data_14,in12_data_13,in12_data_12,in12_data_11,
in12_data_10,in12_data_9,in12_data_8,in12_data_7,in12_data_6,in12_data_5,in12_data_4,gnd,gnd,gnd,gnd,in11_data_15,in11_data_14,in11_data_13,in11_data_12,in11_data_11,in11_data_10,in11_data_9,in11_data_8,in11_data_7,in11_data_6,in11_data_5,in11_data_4,gnd,gnd,gnd,gnd,in10_data_15,
in10_data_14,in10_data_13,in10_data_12,in10_data_11,in10_data_10,in10_data_9,in10_data_8,in10_data_7,in10_data_6,in10_data_5,in10_data_4,gnd,gnd,gnd,gnd,in9_data_15,in9_data_14,in9_data_13,in9_data_12,in9_data_11,in9_data_10,in9_data_9,in9_data_8,in9_data_7,in9_data_6,in9_data_5,
in9_data_4,gnd,gnd,gnd,gnd,in8_data_15,in8_data_14,in8_data_13,in8_data_12,in8_data_11,in8_data_10,in8_data_9,in8_data_8,in8_data_7,in8_data_6,in8_data_5,in8_data_4,gnd,gnd,gnd,gnd,in7_data_15,in7_data_14,in7_data_13,in7_data_12,in7_data_11,in7_data_10,in7_data_9,in7_data_8,in7_data_7,
in7_data_6,in7_data_5,in7_data_4,gnd,gnd,gnd,gnd,in6_data_15,in6_data_14,in6_data_13,in6_data_12,in6_data_11,in6_data_10,in6_data_9,in6_data_8,in6_data_7,in6_data_6,in6_data_5,in6_data_4,gnd,gnd,gnd,gnd,in5_data_15,in5_data_14,in5_data_13,in5_data_12,in5_data_11,in5_data_10,in5_data_9,
in5_data_8,in5_data_7,in5_data_6,in5_data_5,in5_data_4,gnd,gnd,gnd,gnd,in4_data_15,in4_data_14,in4_data_13,in4_data_12,in4_data_11,in4_data_10,in4_data_9,in4_data_8,in4_data_7,in4_data_6,in4_data_5,in4_data_4,gnd,gnd,gnd,gnd,in3_data_15,in3_data_14,in3_data_13,in3_data_12,in3_data_11,
in3_data_10,in3_data_9,in3_data_8,in3_data_7,in3_data_6,in3_data_5,in3_data_4,gnd,gnd,gnd,gnd,in2_data_15,in2_data_14,in2_data_13,in2_data_12,in2_data_11,in2_data_10,in2_data_9,in2_data_8,in2_data_7,in2_data_6,in2_data_5,in2_data_4,gnd,gnd,gnd,gnd,in1_data_15,in1_data_14,in1_data_13,
in1_data_12,in1_data_11,in1_data_10,in1_data_9,in1_data_8,in1_data_7,in1_data_6,in1_data_5,in1_data_4,gnd,gnd,gnd,gnd,in0_data_15,in0_data_14,in0_data_13,in0_data_12,in0_data_11,in0_data_10,in0_data_9,in0_data_8,in0_data_7,in0_data_6,in0_data_5,in0_data_4,gnd,gnd,gnd,gnd}));

endmodule

module CIC_alt_cic_dec_miso (
	state_0,
	dout_1,
	dout_2,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	q_b_170,
	q_b_169,
	q_b_168,
	q_b_167,
	q_b_166,
	q_b_165,
	q_b_164,
	q_b_106,
	q_b_105,
	q_b_104,
	q_b_103,
	q_b_102,
	q_b_101,
	q_b_100,
	q_b_234,
	q_b_233,
	q_b_232,
	q_b_231,
	q_b_230,
	q_b_229,
	q_b_228,
	q_b_42,
	q_b_41,
	q_b_40,
	q_b_39,
	q_b_38,
	q_b_37,
	q_b_36,
	q_b_186,
	q_b_185,
	q_b_184,
	q_b_183,
	q_b_182,
	q_b_181,
	q_b_180,
	q_b_122,
	q_b_121,
	q_b_120,
	q_b_119,
	q_b_118,
	q_b_117,
	q_b_116,
	q_b_250,
	q_b_249,
	q_b_248,
	q_b_247,
	q_b_246,
	q_b_245,
	q_b_244,
	q_b_58,
	q_b_57,
	q_b_56,
	q_b_55,
	q_b_54,
	q_b_53,
	q_b_52,
	q_b_90,
	q_b_89,
	q_b_88,
	q_b_87,
	q_b_86,
	q_b_85,
	q_b_84,
	q_b_154,
	q_b_153,
	q_b_152,
	q_b_151,
	q_b_150,
	q_b_149,
	q_b_148,
	q_b_218,
	q_b_217,
	q_b_216,
	q_b_215,
	q_b_214,
	q_b_213,
	q_b_212,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_74,
	q_b_73,
	q_b_72,
	q_b_71,
	q_b_70,
	q_b_69,
	q_b_68,
	q_b_138,
	q_b_137,
	q_b_136,
	q_b_135,
	q_b_134,
	q_b_133,
	q_b_132,
	q_b_202,
	q_b_201,
	q_b_200,
	q_b_199,
	q_b_198,
	q_b_197,
	q_b_196,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_107,
	q_b_123,
	q_b_91,
	q_b_75,
	q_b_171,
	q_b_187,
	q_b_155,
	q_b_139,
	q_b_235,
	q_b_251,
	q_b_219,
	q_b_203,
	q_b_43,
	q_b_59,
	q_b_27,
	q_b_11,
	q_b_108,
	q_b_172,
	q_b_236,
	q_b_44,
	q_b_124,
	q_b_188,
	q_b_252,
	q_b_60,
	q_b_156,
	q_b_92,
	q_b_220,
	q_b_28,
	q_b_140,
	q_b_76,
	q_b_204,
	q_b_12,
	q_b_173,
	q_b_189,
	q_b_157,
	q_b_141,
	q_b_109,
	q_b_125,
	q_b_93,
	q_b_77,
	q_b_237,
	q_b_253,
	q_b_221,
	q_b_205,
	q_b_45,
	q_b_61,
	q_b_29,
	q_b_13,
	q_b_174,
	q_b_110,
	q_b_238,
	q_b_46,
	q_b_190,
	q_b_126,
	q_b_254,
	q_b_62,
	q_b_94,
	q_b_158,
	q_b_222,
	q_b_30,
	q_b_78,
	q_b_142,
	q_b_206,
	q_b_14,
	q_b_111,
	q_b_127,
	q_b_95,
	q_b_79,
	q_b_175,
	q_b_191,
	q_b_159,
	q_b_143,
	q_b_239,
	q_b_255,
	q_b_223,
	q_b_207,
	q_b_47,
	q_b_63,
	q_b_31,
	q_b_15,
	stall_reg,
	dout_valid,
	channel_out_int_0,
	channel_out_int_1,
	channel_out_int_2,
	channel_out_int_3,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	state_0;
output 	dout_1;
output 	dout_2;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
input 	q_b_170;
input 	q_b_169;
input 	q_b_168;
input 	q_b_167;
input 	q_b_166;
input 	q_b_165;
input 	q_b_164;
input 	q_b_106;
input 	q_b_105;
input 	q_b_104;
input 	q_b_103;
input 	q_b_102;
input 	q_b_101;
input 	q_b_100;
input 	q_b_234;
input 	q_b_233;
input 	q_b_232;
input 	q_b_231;
input 	q_b_230;
input 	q_b_229;
input 	q_b_228;
input 	q_b_42;
input 	q_b_41;
input 	q_b_40;
input 	q_b_39;
input 	q_b_38;
input 	q_b_37;
input 	q_b_36;
input 	q_b_186;
input 	q_b_185;
input 	q_b_184;
input 	q_b_183;
input 	q_b_182;
input 	q_b_181;
input 	q_b_180;
input 	q_b_122;
input 	q_b_121;
input 	q_b_120;
input 	q_b_119;
input 	q_b_118;
input 	q_b_117;
input 	q_b_116;
input 	q_b_250;
input 	q_b_249;
input 	q_b_248;
input 	q_b_247;
input 	q_b_246;
input 	q_b_245;
input 	q_b_244;
input 	q_b_58;
input 	q_b_57;
input 	q_b_56;
input 	q_b_55;
input 	q_b_54;
input 	q_b_53;
input 	q_b_52;
input 	q_b_90;
input 	q_b_89;
input 	q_b_88;
input 	q_b_87;
input 	q_b_86;
input 	q_b_85;
input 	q_b_84;
input 	q_b_154;
input 	q_b_153;
input 	q_b_152;
input 	q_b_151;
input 	q_b_150;
input 	q_b_149;
input 	q_b_148;
input 	q_b_218;
input 	q_b_217;
input 	q_b_216;
input 	q_b_215;
input 	q_b_214;
input 	q_b_213;
input 	q_b_212;
input 	q_b_26;
input 	q_b_25;
input 	q_b_24;
input 	q_b_23;
input 	q_b_22;
input 	q_b_21;
input 	q_b_20;
input 	q_b_74;
input 	q_b_73;
input 	q_b_72;
input 	q_b_71;
input 	q_b_70;
input 	q_b_69;
input 	q_b_68;
input 	q_b_138;
input 	q_b_137;
input 	q_b_136;
input 	q_b_135;
input 	q_b_134;
input 	q_b_133;
input 	q_b_132;
input 	q_b_202;
input 	q_b_201;
input 	q_b_200;
input 	q_b_199;
input 	q_b_198;
input 	q_b_197;
input 	q_b_196;
input 	q_b_10;
input 	q_b_9;
input 	q_b_8;
input 	q_b_7;
input 	q_b_6;
input 	q_b_5;
input 	q_b_4;
input 	q_b_107;
input 	q_b_123;
input 	q_b_91;
input 	q_b_75;
input 	q_b_171;
input 	q_b_187;
input 	q_b_155;
input 	q_b_139;
input 	q_b_235;
input 	q_b_251;
input 	q_b_219;
input 	q_b_203;
input 	q_b_43;
input 	q_b_59;
input 	q_b_27;
input 	q_b_11;
input 	q_b_108;
input 	q_b_172;
input 	q_b_236;
input 	q_b_44;
input 	q_b_124;
input 	q_b_188;
input 	q_b_252;
input 	q_b_60;
input 	q_b_156;
input 	q_b_92;
input 	q_b_220;
input 	q_b_28;
input 	q_b_140;
input 	q_b_76;
input 	q_b_204;
input 	q_b_12;
input 	q_b_173;
input 	q_b_189;
input 	q_b_157;
input 	q_b_141;
input 	q_b_109;
input 	q_b_125;
input 	q_b_93;
input 	q_b_77;
input 	q_b_237;
input 	q_b_253;
input 	q_b_221;
input 	q_b_205;
input 	q_b_45;
input 	q_b_61;
input 	q_b_29;
input 	q_b_13;
input 	q_b_174;
input 	q_b_110;
input 	q_b_238;
input 	q_b_46;
input 	q_b_190;
input 	q_b_126;
input 	q_b_254;
input 	q_b_62;
input 	q_b_94;
input 	q_b_158;
input 	q_b_222;
input 	q_b_30;
input 	q_b_78;
input 	q_b_142;
input 	q_b_206;
input 	q_b_14;
input 	q_b_111;
input 	q_b_127;
input 	q_b_95;
input 	q_b_79;
input 	q_b_175;
input 	q_b_191;
input 	q_b_159;
input 	q_b_143;
input 	q_b_239;
input 	q_b_255;
input 	q_b_223;
input 	q_b_207;
input 	q_b_47;
input 	q_b_63;
input 	q_b_31;
input 	q_b_15;
input 	stall_reg;
output 	dout_valid;
output 	channel_out_int_0;
output 	channel_out_int_1;
output 	channel_out_int_2;
output 	channel_out_int_3;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \ena_sample~q ;
wire \sample_state[0]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[7]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[8]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[9]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ;
wire \fifo_rdreq[10]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[6]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[14]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[2]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[11]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[7]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[3]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[5]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[9]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[13]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[1]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[4]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[8]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[12]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \fifo_rdreq[0]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ;
wire \integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~1 ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~0_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~3 ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~2_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~5 ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~4_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~7 ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~6_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~9 ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~8_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~1 ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~0_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~3 ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~2_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~5 ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~4_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~7 ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~6_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~9 ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~8_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[6]~11_cout ;
wire \Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~1 ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~0_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~3 ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~2_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~5 ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~4_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~7 ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~6_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~9 ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~8_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[6]~11_cout ;
wire \Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~1 ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~0_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~3 ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~2_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~5 ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~4_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~7 ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~6_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~9 ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~8_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[6]~11_cout ;
wire \Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~1 ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~0_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~3 ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~2_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~5 ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~4_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~7 ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~6_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~9 ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~8_combout ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[6]~11_cout ;
wire \Mod0|auto_generated|divider|divider|add_sub_9_result_int[7]~12_combout ;
wire \ena_diff_s[1]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ;
wire \int_channel_cnt_inst|count[1]~q ;
wire \int_channel_cnt_inst|count[0]~q ;
wire \int_channel_cnt_inst|count[2]~q ;
wire \Add1~0_combout ;
wire \int_channel_cnt_inst|count[3]~q ;
wire \Add1~1_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Mux15~6_combout ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \Mux15~9_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \Mux16~7_combout ;
wire \Mux16~8_combout ;
wire \Mux16~9_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \Mux14~6_combout ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \Mux14~9_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Mux13~4_combout ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \Mux13~9_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \Mux12~7_combout ;
wire \Mux12~8_combout ;
wire \Mux12~9_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \Mux11~6_combout ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \Mux11~9_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Mux10~6_combout ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \Mux10~9_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~6_combout ;
wire \Mux9~7_combout ;
wire \Mux9~8_combout ;
wire \Mux9~9_combout ;
wire \Add1~2_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \Mux8~9_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \Mux7~9_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~9_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \Mux5~6_combout ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \Mux5~9_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \Mux4~9_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Mux3~6_combout ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \Mux3~9_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux2~6_combout ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \Mux2~9_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \Mux1~9_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \Mux0~9_combout ;
wire \ena_diff_s~0_combout ;
wire \ena_sample~0_combout ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ;
wire \Equal6~0_combout ;
wire \fifo_rdreq[15]~q ;
wire \Mod0|auto_generated|divider|divider|StageOut[40]~60_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[40]~61_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[39]~62_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[39]~63_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[38]~64_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[38]~65_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[37]~66_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[37]~67_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[36]~68_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[36]~69_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[35]~70_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[35]~71_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[47]~72_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[46]~73_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[45]~74_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[44]~75_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[43]~76_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[43]~77_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[42]~78_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[42]~79_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[54]~80_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[53]~81_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[52]~82_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[51]~83_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[50]~84_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[50]~85_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[49]~86_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[49]~87_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[61]~88_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[60]~89_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[59]~90_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[58]~91_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[57]~92_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[57]~93_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[56]~94_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[56]~95_combout ;
wire \ena_sample~1_combout ;
wire \ena_sample~2_combout ;
wire \ena_sample~3_combout ;
wire \ena_sample~4_combout ;
wire \ena_sample~5_combout ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|Equal0~0_combout ;
wire \ena_sample~6_combout ;
wire \ena_sample~7_combout ;
wire \ena_sample~8_combout ;
wire \ena_sample~9_combout ;
wire \ena_sample~10_combout ;
wire \sample_state~0_combout ;
wire \Equal6~1_combout ;
wire \Equal6~2_combout ;
wire \Equal6~3_combout ;
wire \Equal6~4_combout ;
wire \Equal6~5_combout ;
wire \Equal6~6_combout ;
wire \always5~0_combout ;
wire \Equal6~7_combout ;
wire \Equal6~8_combout ;
wire \Equal6~9_combout ;
wire \Equal6~10_combout ;
wire \Equal6~11_combout ;
wire \Equal6~12_combout ;
wire \Equal6~13_combout ;
wire \Equal6~14_combout ;
wire \Equal6~15_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[54]~96_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[53]~97_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[52]~98_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[61]~99_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[60]~100_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[59]~101_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[47]~102_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[46]~103_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[45]~104_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[44]~105_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[51]~106_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[58]~107_combout ;
wire \latency_cnt[2]~0_combout ;
wire \latency_cnt[0]~3_combout ;
wire \latency_cnt[0]~q ;
wire \latency_cnt[1]~2_combout ;
wire \latency_cnt[1]~q ;
wire \Add2~0_combout ;
wire \latency_cnt[2]~1_combout ;
wire \latency_cnt[2]~q ;
wire \state~0_combout ;
wire \state~1_combout ;
wire \channel_out_int~0_combout ;
wire \channel_out_int[3]~1_combout ;
wire \channel_out_int[3]~2_combout ;
wire \channel_out_int~3_combout ;
wire \Add0~0_combout ;
wire \channel_out_int~4_combout ;
wire \channel_out_int~5_combout ;


CIC_auk_dspip_integrator \integrator[0].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_10(q_b_10),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.stall_reg(stall_reg),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_differentiator \stage_diff[0].auk_dsp_diff (
	.dout_1(dout_1),
	.dout_2(dout_2),
	.dout_3(dout_3),
	.dout_4(dout_4),
	.dout_5(dout_5),
	.dout_6(dout_6),
	.dout_7(dout_7),
	.dout_8(dout_8),
	.dout_9(dout_9),
	.dout_10(dout_10),
	.dout_11(dout_11),
	.dout_12(dout_12),
	.dout_13(dout_13),
	.dout_14(dout_14),
	.dout_15(dout_15),
	.dout_16(dout_16),
	.stall_reg(stall_reg),
	.dout_valid1(dout_valid),
	.ena_diff_s_1(\ena_diff_s[1]~q ),
	.register_fifofifo_data013(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.Mux15(\Mux15~9_combout ),
	.Mux16(\Mux16~9_combout ),
	.Mux14(\Mux14~9_combout ),
	.Mux13(\Mux13~9_combout ),
	.Mux12(\Mux12~9_combout ),
	.Mux11(\Mux11~9_combout ),
	.Mux10(\Mux10~9_combout ),
	.Mux9(\Mux9~9_combout ),
	.Mux8(\Mux8~9_combout ),
	.Mux7(\Mux7~9_combout ),
	.Mux6(\Mux6~9_combout ),
	.Mux5(\Mux5~9_combout ),
	.Mux4(\Mux4~9_combout ),
	.Mux3(\Mux3~9_combout ),
	.Mux2(\Mux2~9_combout ),
	.Mux1(\Mux1~9_combout ),
	.Mux0(\Mux0~9_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_counter_module_33 int_channel_cnt_inst(
	.ena_sample(\ena_sample~q ),
	.stall_reg(stall_reg),
	.count_1(\int_channel_cnt_inst|count[1]~q ),
	.count_0(\int_channel_cnt_inst|count[0]~q ),
	.count_2(\int_channel_cnt_inst|count[2]~q ),
	.count_3(\int_channel_cnt_inst|count[3]~q ),
	.Equal6(\Equal6~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_6 \integrator[15].fifo_regulator (
	.q({\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,
q_unconnected_wire_0}),
	.data({\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.fifo_rdreq_15(\fifo_rdreq[15]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_6 \integrator[15].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[15].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_250(q_b_250),
	.q_b_249(q_b_249),
	.q_b_248(q_b_248),
	.q_b_247(q_b_247),
	.q_b_246(q_b_246),
	.q_b_245(q_b_245),
	.q_b_244(q_b_244),
	.q_b_251(q_b_251),
	.q_b_252(q_b_252),
	.q_b_253(q_b_253),
	.q_b_254(q_b_254),
	.q_b_255(q_b_255),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_5 \integrator[14].fifo_regulator (
	.q({\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_1,q_unconnected_wire_3_1,q_unconnected_wire_2_1,q_unconnected_wire_1_1,
q_unconnected_wire_0_1}),
	.fifo_rdreq_14(\fifo_rdreq[14]~q ),
	.data({\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_5 \integrator[14].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[14].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_234(q_b_234),
	.q_b_233(q_b_233),
	.q_b_232(q_b_232),
	.q_b_231(q_b_231),
	.q_b_230(q_b_230),
	.q_b_229(q_b_229),
	.q_b_228(q_b_228),
	.q_b_235(q_b_235),
	.q_b_236(q_b_236),
	.q_b_237(q_b_237),
	.q_b_238(q_b_238),
	.q_b_239(q_b_239),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_4 \integrator[13].fifo_regulator (
	.q({\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_2,q_unconnected_wire_3_2,q_unconnected_wire_2_2,q_unconnected_wire_1_2,
q_unconnected_wire_0_2}),
	.fifo_rdreq_13(\fifo_rdreq[13]~q ),
	.data({\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_4 \integrator[13].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[13].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_218(q_b_218),
	.q_b_217(q_b_217),
	.q_b_216(q_b_216),
	.q_b_215(q_b_215),
	.q_b_214(q_b_214),
	.q_b_213(q_b_213),
	.q_b_212(q_b_212),
	.q_b_219(q_b_219),
	.q_b_220(q_b_220),
	.q_b_221(q_b_221),
	.q_b_222(q_b_222),
	.q_b_223(q_b_223),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_3 \integrator[12].fifo_regulator (
	.q({\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_3,q_unconnected_wire_3_3,q_unconnected_wire_2_3,q_unconnected_wire_1_3,
q_unconnected_wire_0_3}),
	.fifo_rdreq_12(\fifo_rdreq[12]~q ),
	.data({\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_3 \integrator[12].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[12].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_202(q_b_202),
	.q_b_201(q_b_201),
	.q_b_200(q_b_200),
	.q_b_199(q_b_199),
	.q_b_198(q_b_198),
	.q_b_197(q_b_197),
	.q_b_196(q_b_196),
	.q_b_203(q_b_203),
	.q_b_204(q_b_204),
	.q_b_205(q_b_205),
	.q_b_206(q_b_206),
	.q_b_207(q_b_207),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_2 \integrator[11].fifo_regulator (
	.q({\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_4,q_unconnected_wire_3_4,q_unconnected_wire_2_4,q_unconnected_wire_1_4,
q_unconnected_wire_0_4}),
	.fifo_rdreq_11(\fifo_rdreq[11]~q ),
	.data({\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_2 \integrator[11].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[11].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_186(q_b_186),
	.q_b_185(q_b_185),
	.q_b_184(q_b_184),
	.q_b_183(q_b_183),
	.q_b_182(q_b_182),
	.q_b_181(q_b_181),
	.q_b_180(q_b_180),
	.q_b_187(q_b_187),
	.q_b_188(q_b_188),
	.q_b_189(q_b_189),
	.q_b_190(q_b_190),
	.q_b_191(q_b_191),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_1 \integrator[10].fifo_regulator (
	.q({\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_5,q_unconnected_wire_3_5,q_unconnected_wire_2_5,q_unconnected_wire_1_5,
q_unconnected_wire_0_5}),
	.fifo_rdreq_10(\fifo_rdreq[10]~q ),
	.data({\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_1 \integrator[10].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[10].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_170(q_b_170),
	.q_b_169(q_b_169),
	.q_b_168(q_b_168),
	.q_b_167(q_b_167),
	.q_b_166(q_b_166),
	.q_b_165(q_b_165),
	.q_b_164(q_b_164),
	.q_b_171(q_b_171),
	.q_b_172(q_b_172),
	.q_b_173(q_b_173),
	.q_b_174(q_b_174),
	.q_b_175(q_b_175),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_15 \integrator[9].fifo_regulator (
	.q({\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_6,q_unconnected_wire_3_6,q_unconnected_wire_2_6,q_unconnected_wire_1_6,
q_unconnected_wire_0_6}),
	.fifo_rdreq_9(\fifo_rdreq[9]~q ),
	.data({\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_15 \integrator[9].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[9].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_154(q_b_154),
	.q_b_153(q_b_153),
	.q_b_152(q_b_152),
	.q_b_151(q_b_151),
	.q_b_150(q_b_150),
	.q_b_149(q_b_149),
	.q_b_148(q_b_148),
	.q_b_155(q_b_155),
	.q_b_156(q_b_156),
	.q_b_157(q_b_157),
	.q_b_158(q_b_158),
	.q_b_159(q_b_159),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_14 \integrator[8].fifo_regulator (
	.q({\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_7,q_unconnected_wire_3_7,q_unconnected_wire_2_7,q_unconnected_wire_1_7,
q_unconnected_wire_0_7}),
	.fifo_rdreq_8(\fifo_rdreq[8]~q ),
	.data({\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_14 \integrator[8].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_138(q_b_138),
	.q_b_137(q_b_137),
	.q_b_136(q_b_136),
	.q_b_135(q_b_135),
	.q_b_134(q_b_134),
	.q_b_133(q_b_133),
	.q_b_132(q_b_132),
	.q_b_139(q_b_139),
	.q_b_140(q_b_140),
	.q_b_141(q_b_141),
	.q_b_142(q_b_142),
	.q_b_143(q_b_143),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_13 \integrator[7].fifo_regulator (
	.q({\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_8,q_unconnected_wire_3_8,q_unconnected_wire_2_8,q_unconnected_wire_1_8,
q_unconnected_wire_0_8}),
	.fifo_rdreq_7(\fifo_rdreq[7]~q ),
	.data({\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_13 \integrator[7].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_122(q_b_122),
	.q_b_121(q_b_121),
	.q_b_120(q_b_120),
	.q_b_119(q_b_119),
	.q_b_118(q_b_118),
	.q_b_117(q_b_117),
	.q_b_116(q_b_116),
	.q_b_123(q_b_123),
	.q_b_124(q_b_124),
	.q_b_125(q_b_125),
	.q_b_126(q_b_126),
	.q_b_127(q_b_127),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_12 \integrator[6].fifo_regulator (
	.q({\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_9,q_unconnected_wire_3_9,q_unconnected_wire_2_9,q_unconnected_wire_1_9,
q_unconnected_wire_0_9}),
	.fifo_rdreq_6(\fifo_rdreq[6]~q ),
	.data({\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_12 \integrator[6].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_106(q_b_106),
	.q_b_105(q_b_105),
	.q_b_104(q_b_104),
	.q_b_103(q_b_103),
	.q_b_102(q_b_102),
	.q_b_101(q_b_101),
	.q_b_100(q_b_100),
	.q_b_107(q_b_107),
	.q_b_108(q_b_108),
	.q_b_109(q_b_109),
	.q_b_110(q_b_110),
	.q_b_111(q_b_111),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_11 \integrator[5].fifo_regulator (
	.q({\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_10,q_unconnected_wire_3_10,q_unconnected_wire_2_10,q_unconnected_wire_1_10,
q_unconnected_wire_0_10}),
	.fifo_rdreq_5(\fifo_rdreq[5]~q ),
	.data({\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_11 \integrator[5].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_90(q_b_90),
	.q_b_89(q_b_89),
	.q_b_88(q_b_88),
	.q_b_87(q_b_87),
	.q_b_86(q_b_86),
	.q_b_85(q_b_85),
	.q_b_84(q_b_84),
	.q_b_91(q_b_91),
	.q_b_92(q_b_92),
	.q_b_93(q_b_93),
	.q_b_94(q_b_94),
	.q_b_95(q_b_95),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_10 \integrator[4].fifo_regulator (
	.q({\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_11,q_unconnected_wire_3_11,q_unconnected_wire_2_11,q_unconnected_wire_1_11,
q_unconnected_wire_0_11}),
	.fifo_rdreq_4(\fifo_rdreq[4]~q ),
	.data({\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_10 \integrator[4].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_74(q_b_74),
	.q_b_73(q_b_73),
	.q_b_72(q_b_72),
	.q_b_71(q_b_71),
	.q_b_70(q_b_70),
	.q_b_69(q_b_69),
	.q_b_68(q_b_68),
	.q_b_75(q_b_75),
	.q_b_76(q_b_76),
	.q_b_77(q_b_77),
	.q_b_78(q_b_78),
	.q_b_79(q_b_79),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_9 \integrator[3].fifo_regulator (
	.q({\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_12,q_unconnected_wire_3_12,q_unconnected_wire_2_12,q_unconnected_wire_1_12,
q_unconnected_wire_0_12}),
	.fifo_rdreq_3(\fifo_rdreq[3]~q ),
	.data({\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_9 \integrator[3].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_58(q_b_58),
	.q_b_57(q_b_57),
	.q_b_56(q_b_56),
	.q_b_55(q_b_55),
	.q_b_54(q_b_54),
	.q_b_53(q_b_53),
	.q_b_52(q_b_52),
	.q_b_59(q_b_59),
	.q_b_60(q_b_60),
	.q_b_61(q_b_61),
	.q_b_62(q_b_62),
	.q_b_63(q_b_63),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_8 \integrator[2].fifo_regulator (
	.q({\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_13,q_unconnected_wire_3_13,q_unconnected_wire_2_13,q_unconnected_wire_1_13,
q_unconnected_wire_0_13}),
	.fifo_rdreq_2(\fifo_rdreq[2]~q ),
	.data({\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_8 \integrator[2].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_42(q_b_42),
	.q_b_41(q_b_41),
	.q_b_40(q_b_40),
	.q_b_39(q_b_39),
	.q_b_38(q_b_38),
	.q_b_37(q_b_37),
	.q_b_36(q_b_36),
	.q_b_43(q_b_43),
	.q_b_44(q_b_44),
	.q_b_45(q_b_45),
	.q_b_46(q_b_46),
	.q_b_47(q_b_47),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer_7 \integrator[1].fifo_regulator (
	.q({\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_14,q_unconnected_wire_3_14,q_unconnected_wire_2_14,q_unconnected_wire_1_14,
q_unconnected_wire_0_14}),
	.count_3(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.count_4(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.count_2(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.count_5(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.count_6(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.count_7(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[7]~q ),
	.count_8(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[8]~q ),
	.count_9(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[9]~q ),
	.count_1(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.fifo_rdreq_1(\fifo_rdreq[1]~q ),
	.data({\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.ena_sample(\ena_sample~0_combout ),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_integrator_7 \integrator[1].integrator_inner[0].integration (
	.register_fifofifo_data06(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data05(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data07(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data019(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ),
	.register_fifofifo_data020(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ),
	.register_fifofifo_data021(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ),
	.q_b_26(q_b_26),
	.q_b_25(q_b_25),
	.q_b_24(q_b_24),
	.q_b_23(q_b_23),
	.q_b_22(q_b_22),
	.q_b_21(q_b_21),
	.q_b_20(q_b_20),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_channel_buffer \integrator[0].fifo_regulator (
	.q({\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,q_unconnected_wire_4_15,q_unconnected_wire_3_15,q_unconnected_wire_2_15,q_unconnected_wire_1_15,
q_unconnected_wire_0_15}),
	.fifo_rdreq_0(\fifo_rdreq[0]~q ),
	.data({\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][21]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][20]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][19]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,
\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

CIC_auk_dspip_downsample \integrator[0].j0.vrc_en_0.first_dsample (
	.sample_state_0(\sample_state[0]~q ),
	.count_0(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.count_3(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.count_4(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.count_2(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.count_5(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.count_6(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.count_7(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[7]~q ),
	.count_8(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[8]~q ),
	.count_9(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[9]~q ),
	.count_1(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.stall_reg(stall_reg),
	.ena_sample(\ena_sample~5_combout ),
	.Equal0(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|Equal0~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

dffeas ena_sample(
	.clk(clk),
	.d(\ena_sample~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\ena_sample~q ),
	.prn(vcc));
defparam ena_sample.is_wysiwyg = "true";
defparam ena_sample.power_up = "low";

dffeas \sample_state[0] (
	.clk(clk),
	.d(\sample_state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\sample_state[0]~q ),
	.prn(vcc));
defparam \sample_state[0] .is_wysiwyg = "true";
defparam \sample_state[0] .power_up = "low";

dffeas \fifo_rdreq[10] (
	.clk(clk),
	.d(\Equal6~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[10]~q ),
	.prn(vcc));
defparam \fifo_rdreq[10] .is_wysiwyg = "true";
defparam \fifo_rdreq[10] .power_up = "low";

dffeas \fifo_rdreq[6] (
	.clk(clk),
	.d(\Equal6~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[6]~q ),
	.prn(vcc));
defparam \fifo_rdreq[6] .is_wysiwyg = "true";
defparam \fifo_rdreq[6] .power_up = "low";

dffeas \fifo_rdreq[14] (
	.clk(clk),
	.d(\Equal6~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[14]~q ),
	.prn(vcc));
defparam \fifo_rdreq[14] .is_wysiwyg = "true";
defparam \fifo_rdreq[14] .power_up = "low";

dffeas \fifo_rdreq[2] (
	.clk(clk),
	.d(\Equal6~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[2]~q ),
	.prn(vcc));
defparam \fifo_rdreq[2] .is_wysiwyg = "true";
defparam \fifo_rdreq[2] .power_up = "low";

dffeas \fifo_rdreq[11] (
	.clk(clk),
	.d(\Equal6~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[11]~q ),
	.prn(vcc));
defparam \fifo_rdreq[11] .is_wysiwyg = "true";
defparam \fifo_rdreq[11] .power_up = "low";

dffeas \fifo_rdreq[7] (
	.clk(clk),
	.d(\Equal6~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[7]~q ),
	.prn(vcc));
defparam \fifo_rdreq[7] .is_wysiwyg = "true";
defparam \fifo_rdreq[7] .power_up = "low";

dffeas \fifo_rdreq[3] (
	.clk(clk),
	.d(\Equal6~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[3]~q ),
	.prn(vcc));
defparam \fifo_rdreq[3] .is_wysiwyg = "true";
defparam \fifo_rdreq[3] .power_up = "low";

dffeas \fifo_rdreq[5] (
	.clk(clk),
	.d(\Equal6~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[5]~q ),
	.prn(vcc));
defparam \fifo_rdreq[5] .is_wysiwyg = "true";
defparam \fifo_rdreq[5] .power_up = "low";

dffeas \fifo_rdreq[9] (
	.clk(clk),
	.d(\Equal6~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[9]~q ),
	.prn(vcc));
defparam \fifo_rdreq[9] .is_wysiwyg = "true";
defparam \fifo_rdreq[9] .power_up = "low";

dffeas \fifo_rdreq[13] (
	.clk(clk),
	.d(\Equal6~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[13]~q ),
	.prn(vcc));
defparam \fifo_rdreq[13] .is_wysiwyg = "true";
defparam \fifo_rdreq[13] .power_up = "low";

dffeas \fifo_rdreq[1] (
	.clk(clk),
	.d(\Equal6~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[1]~q ),
	.prn(vcc));
defparam \fifo_rdreq[1] .is_wysiwyg = "true";
defparam \fifo_rdreq[1] .power_up = "low";

dffeas \fifo_rdreq[4] (
	.clk(clk),
	.d(\Equal6~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[4]~q ),
	.prn(vcc));
defparam \fifo_rdreq[4] .is_wysiwyg = "true";
defparam \fifo_rdreq[4] .power_up = "low";

dffeas \fifo_rdreq[8] (
	.clk(clk),
	.d(\Equal6~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[8]~q ),
	.prn(vcc));
defparam \fifo_rdreq[8] .is_wysiwyg = "true";
defparam \fifo_rdreq[8] .power_up = "low";

dffeas \fifo_rdreq[12] (
	.clk(clk),
	.d(\Equal6~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[12]~q ),
	.prn(vcc));
defparam \fifo_rdreq[12] .is_wysiwyg = "true";
defparam \fifo_rdreq[12] .power_up = "low";

dffeas \fifo_rdreq[0] (
	.clk(clk),
	.d(\Equal6~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\ena_sample~q ),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[0]~q ),
	.prn(vcc));
defparam \fifo_rdreq[0] .is_wysiwyg = "true";
defparam \fifo_rdreq[0] .power_up = "low";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~0 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~1 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~0 .lut_mask = 16'h55AA;
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~2 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~1 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~3 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~2 .lut_mask = 16'h5A5F;
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~4 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~3 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~5 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~4 .lut_mask = 16'h5AAF;
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~6 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~5 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~6_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~7 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~6 .lut_mask = 16'h5A5F;
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~8 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~7 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~8_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~9 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~8 .lut_mask = 16'h5AAF;
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~9 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10 .lut_mask = 16'h0F0F;
defparam \Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~0 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[35]~70_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[35]~71_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~1 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~0 .lut_mask = 16'h77EE;
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[36]~68_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[36]~69_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~1 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~3 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[37]~66_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[37]~67_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~3 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~5 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~6 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[38]~64_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[38]~65_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~5 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~6_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~7 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~6 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~8 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[39]~62_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[39]~63_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~7 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~8_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~9 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~8 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_6_result_int[6]~11 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[40]~60_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[40]~61_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~9 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[6]~11_cout ));
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[6]~11 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[6]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[6]~11_cout ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~0 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[42]~78_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[42]~79_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~1 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~0 .lut_mask = 16'h77EE;
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[43]~76_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[43]~77_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~1 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~3 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[44]~105_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[44]~75_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~3 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~5 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~6 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[45]~104_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[45]~74_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~5 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~6_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~7 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~6 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~8 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[46]~103_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[46]~73_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~7 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~8_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~9 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~8 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_7_result_int[6]~11 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[47]~102_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[47]~72_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~9 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[6]~11_cout ));
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[6]~11 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[6]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[6]~11_cout ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~0 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[49]~86_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[49]~87_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~1 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~0 .lut_mask = 16'h77EE;
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[50]~84_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[50]~85_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~1 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~3 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[51]~106_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[51]~83_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~3 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~5 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~6 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[52]~98_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[52]~82_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~5 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~6_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~7 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~6 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~8 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[53]~97_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[53]~81_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~7 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~8_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~9 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~8 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_8_result_int[6]~11 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[54]~96_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[54]~80_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~9 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[6]~11_cout ));
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[6]~11 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[6]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[6]~11_cout ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~0 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[56]~94_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[56]~95_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~1 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~0 .lut_mask = 16'h77EE;
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[57]~92_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[57]~93_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~1 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~3 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[58]~107_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[58]~91_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~3 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~5 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~6 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[59]~101_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[59]~90_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~5 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~6_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~7 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~6 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~8 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[60]~100_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[60]~89_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~7 ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~8_combout ),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~9 ));
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~8 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_9_result_int[6]~11 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[61]~99_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[61]~88_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~9 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[6]~11_cout ));
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[6]~11 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[6]~11 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|add_sub_9_result_int[7]~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[6]~11_cout ),
	.combout(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[7]~12_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[7]~12 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|add_sub_9_result_int[7]~12 .sum_lutc_input = "cin";

dffeas \ena_diff_s[1] (
	.clk(clk),
	.d(\ena_diff_s~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~1_combout ),
	.q(\ena_diff_s[1]~q ),
	.prn(vcc));
defparam \ena_diff_s[1] .is_wysiwyg = "true";
defparam \ena_diff_s[1] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(\int_channel_cnt_inst|count[1]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[2]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'hC33C;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\int_channel_cnt_inst|count[2]~q ),
	.datab(\int_channel_cnt_inst|count[1]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[3]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~0 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hFFDE;
defparam \Mux15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~1 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux15~0_combout ),
	.datad(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
defparam \Mux15~1 .lut_mask = 16'hFFBE;
defparam \Mux15~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~2 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
defparam \Mux15~2 .lut_mask = 16'hFFDE;
defparam \Mux15~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~3 (
	.dataa(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux15~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
defparam \Mux15~3 .lut_mask = 16'hFFBE;
defparam \Mux15~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~4 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
defparam \Mux15~4 .lut_mask = 16'hFFDE;
defparam \Mux15~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~5 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux15~4_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
defparam \Mux15~5 .lut_mask = 16'hFFBE;
defparam \Mux15~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mux15~3_combout ),
	.datac(\Mux15~5_combout ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
defparam \Mux15~6 .lut_mask = 16'hFDFE;
defparam \Mux15~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~7 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
defparam \Mux15~7 .lut_mask = 16'hFFDE;
defparam \Mux15~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~8 (
	.dataa(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux15~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
defparam \Mux15~8 .lut_mask = 16'hFFBE;
defparam \Mux15~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux15~9 (
	.dataa(\Mux15~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux15~6_combout ),
	.datad(\Mux15~8_combout ),
	.cin(gnd),
	.combout(\Mux15~9_combout ),
	.cout());
defparam \Mux15~9 .lut_mask = 16'hFFBE;
defparam \Mux15~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~0 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'hFDFE;
defparam \Mux16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~1 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux16~0_combout ),
	.datad(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
defparam \Mux16~1 .lut_mask = 16'hFFBE;
defparam \Mux16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~2 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
defparam \Mux16~2 .lut_mask = 16'hFDFE;
defparam \Mux16~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~3 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux16~2_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
defparam \Mux16~3 .lut_mask = 16'hFFBE;
defparam \Mux16~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~4 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
defparam \Mux16~4 .lut_mask = 16'hFDFE;
defparam \Mux16~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~5 (
	.dataa(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux16~4_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
defparam \Mux16~5 .lut_mask = 16'hFFBE;
defparam \Mux16~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~6 (
	.dataa(\Add1~0_combout ),
	.datab(\Mux16~3_combout ),
	.datac(\Add1~1_combout ),
	.datad(\Mux16~5_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
defparam \Mux16~6 .lut_mask = 16'hFFDE;
defparam \Mux16~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~7 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
defparam \Mux16~7 .lut_mask = 16'hFDFE;
defparam \Mux16~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux16~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
defparam \Mux16~8 .lut_mask = 16'hFFBE;
defparam \Mux16~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~9 (
	.dataa(\Mux16~1_combout ),
	.datab(\Add1~0_combout ),
	.datac(\Mux16~6_combout ),
	.datad(\Mux16~8_combout ),
	.cin(gnd),
	.combout(\Mux16~9_combout ),
	.cout());
defparam \Mux16~9 .lut_mask = 16'hFFBE;
defparam \Mux16~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~0 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
defparam \Mux14~0 .lut_mask = 16'hFDFE;
defparam \Mux14~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~1 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux14~0_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
defparam \Mux14~1 .lut_mask = 16'hFFBE;
defparam \Mux14~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~2 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
defparam \Mux14~2 .lut_mask = 16'hFDFE;
defparam \Mux14~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~3 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux14~2_combout ),
	.datad(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
defparam \Mux14~3 .lut_mask = 16'hFFBE;
defparam \Mux14~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~4 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
defparam \Mux14~4 .lut_mask = 16'hFDFE;
defparam \Mux14~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~5 (
	.dataa(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux14~4_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
defparam \Mux14~5 .lut_mask = 16'hFFBE;
defparam \Mux14~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~6 (
	.dataa(\Add1~1_combout ),
	.datab(\Mux14~3_combout ),
	.datac(\Add1~0_combout ),
	.datad(\Mux14~5_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
defparam \Mux14~6 .lut_mask = 16'hFFDE;
defparam \Mux14~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~7 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
defparam \Mux14~7 .lut_mask = 16'hFDFE;
defparam \Mux14~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux14~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
defparam \Mux14~8 .lut_mask = 16'hFFBE;
defparam \Mux14~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux14~9 (
	.dataa(\Mux14~1_combout ),
	.datab(\Add1~1_combout ),
	.datac(\Mux14~6_combout ),
	.datad(\Mux14~8_combout ),
	.cin(gnd),
	.combout(\Mux14~9_combout ),
	.cout());
defparam \Mux14~9 .lut_mask = 16'hFFBE;
defparam \Mux14~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~0 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hFFDE;
defparam \Mux13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~1 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux13~0_combout ),
	.datad(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
defparam \Mux13~1 .lut_mask = 16'hFFBE;
defparam \Mux13~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~2 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
defparam \Mux13~2 .lut_mask = 16'hFFDE;
defparam \Mux13~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~3 (
	.dataa(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux13~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
defparam \Mux13~3 .lut_mask = 16'hFFBE;
defparam \Mux13~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~4 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
defparam \Mux13~4 .lut_mask = 16'hFFDE;
defparam \Mux13~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~5 (
	.dataa(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux13~4_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
defparam \Mux13~5 .lut_mask = 16'hFFBE;
defparam \Mux13~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mux13~3_combout ),
	.datac(\Mux13~5_combout ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
defparam \Mux13~6 .lut_mask = 16'hFDFE;
defparam \Mux13~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~7 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
defparam \Mux13~7 .lut_mask = 16'hFFDE;
defparam \Mux13~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~8 (
	.dataa(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux13~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
defparam \Mux13~8 .lut_mask = 16'hFFBE;
defparam \Mux13~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux13~9 (
	.dataa(\Mux13~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux13~6_combout ),
	.datad(\Mux13~8_combout ),
	.cin(gnd),
	.combout(\Mux13~9_combout ),
	.cout());
defparam \Mux13~9 .lut_mask = 16'hFFBE;
defparam \Mux13~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~0 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hFDFE;
defparam \Mux12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~1 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux12~0_combout ),
	.datad(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
defparam \Mux12~1 .lut_mask = 16'hFFBE;
defparam \Mux12~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~2 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
defparam \Mux12~2 .lut_mask = 16'hFDFE;
defparam \Mux12~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~3 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux12~2_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
defparam \Mux12~3 .lut_mask = 16'hFFBE;
defparam \Mux12~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~4 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
defparam \Mux12~4 .lut_mask = 16'hFDFE;
defparam \Mux12~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~5 (
	.dataa(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux12~4_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
defparam \Mux12~5 .lut_mask = 16'hFFBE;
defparam \Mux12~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~6 (
	.dataa(\Add1~0_combout ),
	.datab(\Mux12~3_combout ),
	.datac(\Add1~1_combout ),
	.datad(\Mux12~5_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
defparam \Mux12~6 .lut_mask = 16'hFFDE;
defparam \Mux12~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~7 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
defparam \Mux12~7 .lut_mask = 16'hFDFE;
defparam \Mux12~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux12~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
defparam \Mux12~8 .lut_mask = 16'hFFBE;
defparam \Mux12~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux12~9 (
	.dataa(\Mux12~1_combout ),
	.datab(\Add1~0_combout ),
	.datac(\Mux12~6_combout ),
	.datad(\Mux12~8_combout ),
	.cin(gnd),
	.combout(\Mux12~9_combout ),
	.cout());
defparam \Mux12~9 .lut_mask = 16'hFFBE;
defparam \Mux12~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~0 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hFFDE;
defparam \Mux11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~1 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux11~0_combout ),
	.datad(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
defparam \Mux11~1 .lut_mask = 16'hFFBE;
defparam \Mux11~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~2 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
defparam \Mux11~2 .lut_mask = 16'hFFDE;
defparam \Mux11~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~3 (
	.dataa(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux11~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
defparam \Mux11~3 .lut_mask = 16'hFFBE;
defparam \Mux11~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~4 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
defparam \Mux11~4 .lut_mask = 16'hFFDE;
defparam \Mux11~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~5 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux11~4_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
defparam \Mux11~5 .lut_mask = 16'hFFBE;
defparam \Mux11~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mux11~3_combout ),
	.datac(\Mux11~5_combout ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
defparam \Mux11~6 .lut_mask = 16'hFDFE;
defparam \Mux11~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~7 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
defparam \Mux11~7 .lut_mask = 16'hFFDE;
defparam \Mux11~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~8 (
	.dataa(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux11~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
defparam \Mux11~8 .lut_mask = 16'hFFBE;
defparam \Mux11~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux11~9 (
	.dataa(\Mux11~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux11~6_combout ),
	.datad(\Mux11~8_combout ),
	.cin(gnd),
	.combout(\Mux11~9_combout ),
	.cout());
defparam \Mux11~9 .lut_mask = 16'hFFBE;
defparam \Mux11~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~0 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hFDFE;
defparam \Mux10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~1 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux10~0_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
defparam \Mux10~1 .lut_mask = 16'hFFBE;
defparam \Mux10~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~2 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
defparam \Mux10~2 .lut_mask = 16'hFDFE;
defparam \Mux10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~3 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux10~2_combout ),
	.datad(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
defparam \Mux10~3 .lut_mask = 16'hFFBE;
defparam \Mux10~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~4 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
defparam \Mux10~4 .lut_mask = 16'hFDFE;
defparam \Mux10~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~5 (
	.dataa(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux10~4_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
defparam \Mux10~5 .lut_mask = 16'hFFBE;
defparam \Mux10~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~6 (
	.dataa(\Add1~1_combout ),
	.datab(\Mux10~3_combout ),
	.datac(\Add1~0_combout ),
	.datad(\Mux10~5_combout ),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
defparam \Mux10~6 .lut_mask = 16'hFFDE;
defparam \Mux10~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~7 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
defparam \Mux10~7 .lut_mask = 16'hFDFE;
defparam \Mux10~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux10~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
defparam \Mux10~8 .lut_mask = 16'hFFBE;
defparam \Mux10~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux10~9 (
	.dataa(\Mux10~1_combout ),
	.datab(\Add1~1_combout ),
	.datac(\Mux10~6_combout ),
	.datad(\Mux10~8_combout ),
	.cin(gnd),
	.combout(\Mux10~9_combout ),
	.cout());
defparam \Mux10~9 .lut_mask = 16'hFFBE;
defparam \Mux10~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~0 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hFFDE;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~1 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux9~0_combout ),
	.datad(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
defparam \Mux9~1 .lut_mask = 16'hFFBE;
defparam \Mux9~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~2 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
defparam \Mux9~2 .lut_mask = 16'hFFDE;
defparam \Mux9~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~3 (
	.dataa(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux9~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
defparam \Mux9~3 .lut_mask = 16'hFFBE;
defparam \Mux9~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~4 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
defparam \Mux9~4 .lut_mask = 16'hFFDE;
defparam \Mux9~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~5 (
	.dataa(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux9~4_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
defparam \Mux9~5 .lut_mask = 16'hFFBE;
defparam \Mux9~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mux9~3_combout ),
	.datac(\Mux9~5_combout ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
defparam \Mux9~6 .lut_mask = 16'hFDFE;
defparam \Mux9~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~7 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
defparam \Mux9~7 .lut_mask = 16'hFFDE;
defparam \Mux9~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~8 (
	.dataa(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux9~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
defparam \Mux9~8 .lut_mask = 16'hFFBE;
defparam \Mux9~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~9 (
	.dataa(\Mux9~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux9~6_combout ),
	.datad(\Mux9~8_combout ),
	.cin(gnd),
	.combout(\Mux9~9_combout ),
	.cout());
defparam \Mux9~9 .lut_mask = 16'hFFBE;
defparam \Mux9~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\int_channel_cnt_inst|count[1]~q ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~0 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hFFDE;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~1 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux8~0_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
defparam \Mux8~1 .lut_mask = 16'hFFBE;
defparam \Mux8~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~2 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
defparam \Mux8~2 .lut_mask = 16'hFFDE;
defparam \Mux8~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~3 (
	.dataa(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux8~2_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
defparam \Mux8~3 .lut_mask = 16'hFFBE;
defparam \Mux8~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~4 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
defparam \Mux8~4 .lut_mask = 16'hFFDE;
defparam \Mux8~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~5 (
	.dataa(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux8~4_combout ),
	.datad(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
defparam \Mux8~5 .lut_mask = 16'hFFBE;
defparam \Mux8~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~6 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mux8~3_combout ),
	.datac(\Add1~0_combout ),
	.datad(\Mux8~5_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
defparam \Mux8~6 .lut_mask = 16'hFFDE;
defparam \Mux8~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~7 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
defparam \Mux8~7 .lut_mask = 16'hFFDE;
defparam \Mux8~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux8~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
defparam \Mux8~8 .lut_mask = 16'hFFBE;
defparam \Mux8~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux8~9 (
	.dataa(\Mux8~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux8~6_combout ),
	.datad(\Mux8~8_combout ),
	.cin(gnd),
	.combout(\Mux8~9_combout ),
	.cout());
defparam \Mux8~9 .lut_mask = 16'hFFBE;
defparam \Mux8~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hFFDE;
defparam \Mux7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~1 (
	.dataa(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux7~0_combout ),
	.datad(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hFFBE;
defparam \Mux7~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~2 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
defparam \Mux7~2 .lut_mask = 16'hFFDE;
defparam \Mux7~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~3 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux7~2_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
defparam \Mux7~3 .lut_mask = 16'hFFBE;
defparam \Mux7~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~4 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
defparam \Mux7~4 .lut_mask = 16'hFFDE;
defparam \Mux7~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~5 (
	.dataa(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux7~4_combout ),
	.datad(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
defparam \Mux7~5 .lut_mask = 16'hFFBE;
defparam \Mux7~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~6 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mux7~3_combout ),
	.datac(\Add1~1_combout ),
	.datad(\Mux7~5_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
defparam \Mux7~6 .lut_mask = 16'hFFDE;
defparam \Mux7~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~7 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
defparam \Mux7~7 .lut_mask = 16'hFFDE;
defparam \Mux7~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~8 (
	.dataa(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux7~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
defparam \Mux7~8 .lut_mask = 16'hFFBE;
defparam \Mux7~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux7~9 (
	.dataa(\Mux7~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux7~6_combout ),
	.datad(\Mux7~8_combout ),
	.cin(gnd),
	.combout(\Mux7~9_combout ),
	.cout());
defparam \Mux7~9 .lut_mask = 16'hFFBE;
defparam \Mux7~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hFFDE;
defparam \Mux6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~1 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux6~0_combout ),
	.datad(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hFFBE;
defparam \Mux6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~2 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hFFDE;
defparam \Mux6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~3 (
	.dataa(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux6~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
defparam \Mux6~3 .lut_mask = 16'hFFBE;
defparam \Mux6~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~4 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
defparam \Mux6~4 .lut_mask = 16'hFFDE;
defparam \Mux6~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~5 (
	.dataa(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux6~4_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
defparam \Mux6~5 .lut_mask = 16'hFFBE;
defparam \Mux6~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mux6~3_combout ),
	.datac(\Mux6~5_combout ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
defparam \Mux6~6 .lut_mask = 16'hFDFE;
defparam \Mux6~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~7 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
defparam \Mux6~7 .lut_mask = 16'hFFDE;
defparam \Mux6~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~8 (
	.dataa(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux6~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
defparam \Mux6~8 .lut_mask = 16'hFFBE;
defparam \Mux6~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux6~9 (
	.dataa(\Mux6~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux6~6_combout ),
	.datad(\Mux6~8_combout ),
	.cin(gnd),
	.combout(\Mux6~9_combout ),
	.cout());
defparam \Mux6~9 .lut_mask = 16'hFFBE;
defparam \Mux6~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hFFDE;
defparam \Mux5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux5~0_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFFBE;
defparam \Mux5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~2 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
defparam \Mux5~2 .lut_mask = 16'hFFDE;
defparam \Mux5~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~3 (
	.dataa(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux5~2_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
defparam \Mux5~3 .lut_mask = 16'hFFBE;
defparam \Mux5~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~4 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
defparam \Mux5~4 .lut_mask = 16'hFFDE;
defparam \Mux5~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~5 (
	.dataa(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux5~4_combout ),
	.datad(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
defparam \Mux5~5 .lut_mask = 16'hFFBE;
defparam \Mux5~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~6 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mux5~3_combout ),
	.datac(\Add1~0_combout ),
	.datad(\Mux5~5_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
defparam \Mux5~6 .lut_mask = 16'hFFDE;
defparam \Mux5~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~7 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
defparam \Mux5~7 .lut_mask = 16'hFFDE;
defparam \Mux5~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux5~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
defparam \Mux5~8 .lut_mask = 16'hFFBE;
defparam \Mux5~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux5~9 (
	.dataa(\Mux5~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux5~6_combout ),
	.datad(\Mux5~8_combout ),
	.cin(gnd),
	.combout(\Mux5~9_combout ),
	.cout());
defparam \Mux5~9 .lut_mask = 16'hFFBE;
defparam \Mux5~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hFFDE;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux4~0_combout ),
	.datad(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hFFBE;
defparam \Mux4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~2 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
defparam \Mux4~2 .lut_mask = 16'hFFDE;
defparam \Mux4~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~3 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux4~2_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
defparam \Mux4~3 .lut_mask = 16'hFFBE;
defparam \Mux4~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~4 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
defparam \Mux4~4 .lut_mask = 16'hFFDE;
defparam \Mux4~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~5 (
	.dataa(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux4~4_combout ),
	.datad(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
defparam \Mux4~5 .lut_mask = 16'hFFBE;
defparam \Mux4~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~6 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mux4~3_combout ),
	.datac(\Add1~1_combout ),
	.datad(\Mux4~5_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
defparam \Mux4~6 .lut_mask = 16'hFFDE;
defparam \Mux4~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~7 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
defparam \Mux4~7 .lut_mask = 16'hFFDE;
defparam \Mux4~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~8 (
	.dataa(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux4~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
defparam \Mux4~8 .lut_mask = 16'hFFBE;
defparam \Mux4~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux4~9 (
	.dataa(\Mux4~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux4~6_combout ),
	.datad(\Mux4~8_combout ),
	.cin(gnd),
	.combout(\Mux4~9_combout ),
	.cout());
defparam \Mux4~9 .lut_mask = 16'hFFBE;
defparam \Mux4~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFFDE;
defparam \Mux3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux3~0_combout ),
	.datad(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hFFBE;
defparam \Mux3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~2 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
defparam \Mux3~2 .lut_mask = 16'hFFDE;
defparam \Mux3~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~3 (
	.dataa(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux3~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
defparam \Mux3~3 .lut_mask = 16'hFFBE;
defparam \Mux3~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~4 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
defparam \Mux3~4 .lut_mask = 16'hFFDE;
defparam \Mux3~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~5 (
	.dataa(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux3~4_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
defparam \Mux3~5 .lut_mask = 16'hFFBE;
defparam \Mux3~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mux3~3_combout ),
	.datac(\Mux3~5_combout ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
defparam \Mux3~6 .lut_mask = 16'hFDFE;
defparam \Mux3~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~7 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
defparam \Mux3~7 .lut_mask = 16'hFFDE;
defparam \Mux3~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~8 (
	.dataa(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux3~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
defparam \Mux3~8 .lut_mask = 16'hFFBE;
defparam \Mux3~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux3~9 (
	.dataa(\Mux3~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux3~6_combout ),
	.datad(\Mux3~8_combout ),
	.cin(gnd),
	.combout(\Mux3~9_combout ),
	.cout());
defparam \Mux3~9 .lut_mask = 16'hFFBE;
defparam \Mux3~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFFDE;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux2~0_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hFFBE;
defparam \Mux2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~2 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hFFDE;
defparam \Mux2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~3 (
	.dataa(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux2~2_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
defparam \Mux2~3 .lut_mask = 16'hFFBE;
defparam \Mux2~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~4 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
defparam \Mux2~4 .lut_mask = 16'hFFDE;
defparam \Mux2~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~5 (
	.dataa(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux2~4_combout ),
	.datad(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
defparam \Mux2~5 .lut_mask = 16'hFFBE;
defparam \Mux2~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~6 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mux2~3_combout ),
	.datac(\Add1~0_combout ),
	.datad(\Mux2~5_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
defparam \Mux2~6 .lut_mask = 16'hFFDE;
defparam \Mux2~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~7 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datac(\Add1~2_combout ),
	.datad(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
defparam \Mux2~7 .lut_mask = 16'hFFDE;
defparam \Mux2~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux2~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
defparam \Mux2~8 .lut_mask = 16'hFFBE;
defparam \Mux2~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~9 (
	.dataa(\Mux2~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux2~6_combout ),
	.datad(\Mux2~8_combout ),
	.cin(gnd),
	.combout(\Mux2~9_combout ),
	.cout());
defparam \Mux2~9 .lut_mask = 16'hFFBE;
defparam \Mux2~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux1~0_combout ),
	.datad(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~2 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hFFDE;
defparam \Mux1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~3 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux1~2_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
defparam \Mux1~3 .lut_mask = 16'hFFBE;
defparam \Mux1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~4 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
defparam \Mux1~4 .lut_mask = 16'hFFDE;
defparam \Mux1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~5 (
	.dataa(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux1~4_combout ),
	.datad(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
defparam \Mux1~5 .lut_mask = 16'hFFBE;
defparam \Mux1~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~6 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mux1~3_combout ),
	.datac(\Add1~1_combout ),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
defparam \Mux1~6 .lut_mask = 16'hFFDE;
defparam \Mux1~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~7 (
	.dataa(\Add1~2_combout ),
	.datab(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
defparam \Mux1~7 .lut_mask = 16'hFFDE;
defparam \Mux1~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~8 (
	.dataa(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.datab(\Add1~2_combout ),
	.datac(\Mux1~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
defparam \Mux1~8 .lut_mask = 16'hFFBE;
defparam \Mux1~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux1~9 (
	.dataa(\Mux1~1_combout ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(\Mux1~6_combout ),
	.datad(\Mux1~8_combout ),
	.cin(gnd),
	.combout(\Mux1~9_combout ),
	.cout());
defparam \Mux1~9 .lut_mask = 16'hFFBE;
defparam \Mux1~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[13].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\integrator[9].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux0~0_combout ),
	.datad(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[11].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[15].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFFDE;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux0~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hFFBE;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~4 (
	.dataa(\Add1~1_combout ),
	.datab(\integrator[10].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datac(\Add1~0_combout ),
	.datad(\integrator[14].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'hFFDE;
defparam \Mux0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~5 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datab(\Add1~1_combout ),
	.datac(\Mux0~4_combout ),
	.datad(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
defparam \Mux0~5 .lut_mask = 16'hFFBE;
defparam \Mux0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mux0~3_combout ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\Mux0~5_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
defparam \Mux0~6 .lut_mask = 16'hFFFD;
defparam \Mux0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~7 (
	.dataa(\Add1~0_combout ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datac(\Add1~1_combout ),
	.datad(\integrator[12].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
defparam \Mux0~7 .lut_mask = 16'hFFDE;
defparam \Mux0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~8 (
	.dataa(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.datab(\Add1~0_combout ),
	.datac(\Mux0~7_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
defparam \Mux0~8 .lut_mask = 16'hFFBE;
defparam \Mux0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~9 (
	.dataa(\Mux0~1_combout ),
	.datab(\Add1~2_combout ),
	.datac(\Mux0~6_combout ),
	.datad(\Mux0~8_combout ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
defparam \Mux0~9 .lut_mask = 16'hFFBE;
defparam \Mux0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_diff_s~0 (
	.dataa(reset_n),
	.datab(\ena_sample~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ena_diff_s~0_combout ),
	.cout());
defparam \ena_diff_s~0 .lut_mask = 16'hEEEE;
defparam \ena_diff_s~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~0 (
	.dataa(\sample_state[0]~q ),
	.datab(gnd),
	.datac(stall_reg),
	.datad(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.cin(gnd),
	.combout(\ena_sample~0_combout ),
	.cout());
defparam \ena_sample~0 .lut_mask = 16'hAFFF;
defparam \ena_sample~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~0 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
defparam \Equal6~0 .lut_mask = 16'hFFFE;
defparam \Equal6~0 .sum_lutc_input = "datac";

dffeas \fifo_rdreq[15] (
	.clk(clk),
	.d(\always5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[15]~q ),
	.prn(vcc));
defparam \fifo_rdreq[15] .is_wysiwyg = "true";
defparam \fifo_rdreq[15] .power_up = "low";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[40]~60 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[9]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[40]~60_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[40]~60 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[40]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[40]~61 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[5]~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[40]~61_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[40]~61 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[40]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[39]~62 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[8]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[39]~62_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[39]~62 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[39]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[39]~63 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[39]~63_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[39]~63 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[39]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[38]~64 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[7]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[38]~64_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[38]~64 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[38]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[38]~65 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[38]~65_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[38]~65 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[38]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[37]~66 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[37]~66_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[37]~66 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[37]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[37]~67 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[37]~67_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[37]~67 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[37]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[36]~68 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[36]~68_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[36]~68 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[36]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[36]~69 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[36]~69_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[36]~69 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[36]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[35]~70 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[35]~70_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[35]~70 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[35]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[35]~71 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[35]~71_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[35]~71 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[35]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[47]~72 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[5]~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[47]~72_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[47]~72 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[47]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[46]~73 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[46]~73_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[46]~73 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[46]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[45]~74 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[45]~74_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[45]~74 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[45]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[44]~75 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[44]~75_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[44]~75 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[44]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[43]~76 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[43]~76_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[43]~76 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[43]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[43]~77 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[43]~77_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[43]~77 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[43]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[42]~78 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[42]~78_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[42]~78 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[42]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[42]~79 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[42]~79_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[42]~79 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[42]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[54]~80 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[5]~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[54]~80_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[54]~80 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[54]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[53]~81 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[53]~81_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[53]~81 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[53]~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[52]~82 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[52]~82_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[52]~82 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[52]~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[51]~83 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[51]~83_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[51]~83 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[51]~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[50]~84 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[50]~84_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[50]~84 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[50]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[50]~85 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[50]~85_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[50]~85 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[50]~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[49]~86 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[49]~86_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[49]~86 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[49]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[49]~87 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[49]~87_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[49]~87 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[49]~87 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[61]~88 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[5]~8_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[61]~88_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[61]~88 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[61]~88 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[60]~89 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[60]~89_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[60]~89 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[60]~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[59]~90 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[59]~90_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[59]~90 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[59]~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[58]~91 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[58]~91_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[58]~91 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[58]~91 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[57]~92 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[57]~92_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[57]~92 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[57]~92 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[57]~93 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[57]~93_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[57]~93 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[57]~93 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[56]~94 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[56]~94_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[56]~94 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[56]~94 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[56]~95 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[56]~95_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[56]~95 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[56]~95 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~1 (
	.dataa(\ena_sample~q ),
	.datab(stall_reg),
	.datac(gnd),
	.datad(\sample_state[0]~q ),
	.cin(gnd),
	.combout(\ena_sample~1_combout ),
	.cout());
defparam \ena_sample~1 .lut_mask = 16'hEEFF;
defparam \ena_sample~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~2 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[3]~4_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[4]~6_combout ),
	.datad(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.cin(gnd),
	.combout(\ena_sample~2_combout ),
	.cout());
defparam \ena_sample~2 .lut_mask = 16'h27FF;
defparam \ena_sample~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~3 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[1]~0_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[2]~2_combout ),
	.datad(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.cin(gnd),
	.combout(\ena_sample~3_combout ),
	.cout());
defparam \ena_sample~3 .lut_mask = 16'hBFFF;
defparam \ena_sample~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[60]~100_combout ),
	.datab(\ena_sample~3_combout ),
	.datac(\Mod0|auto_generated|divider|divider|StageOut[59]~101_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[58]~107_combout ),
	.cin(gnd),
	.combout(\ena_sample~4_combout ),
	.cout());
defparam \ena_sample~4 .lut_mask = 16'hDFFF;
defparam \ena_sample~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datad(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.cin(gnd),
	.combout(\ena_sample~5_combout ),
	.cout());
defparam \ena_sample~5 .lut_mask = 16'h0FFF;
defparam \ena_sample~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~6 (
	.dataa(\ena_sample~5_combout ),
	.datab(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[9]~q ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|Equal0~0_combout ),
	.datad(\ena_sample~0_combout ),
	.cin(gnd),
	.combout(\ena_sample~6_combout ),
	.cout());
defparam \ena_sample~6 .lut_mask = 16'hFFBF;
defparam \ena_sample~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~7 (
	.dataa(\ena_sample~2_combout ),
	.datab(\ena_sample~4_combout ),
	.datac(\ena_sample~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ena_sample~7_combout ),
	.cout());
defparam \ena_sample~7 .lut_mask = 16'hFEFE;
defparam \ena_sample~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~8 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[1]~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[2]~2_combout ),
	.datac(\ena_sample~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ena_sample~8_combout ),
	.cout());
defparam \ena_sample~8 .lut_mask = 16'hF7F7;
defparam \ena_sample~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~9 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[3]~4_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[4]~6_combout ),
	.datac(\ena_sample~8_combout ),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[5]~8_combout ),
	.cin(gnd),
	.combout(\ena_sample~9_combout ),
	.cout());
defparam \ena_sample~9 .lut_mask = 16'hF7FF;
defparam \ena_sample~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ena_sample~10 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_9_result_int[7]~12_combout ),
	.datab(\ena_sample~1_combout ),
	.datac(\ena_sample~7_combout ),
	.datad(\ena_sample~9_combout ),
	.cin(gnd),
	.combout(\ena_sample~10_combout ),
	.cout());
defparam \ena_sample~10 .lut_mask = 16'hFFD8;
defparam \ena_sample~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sample_state~0 (
	.dataa(\sample_state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\sample_state~0_combout ),
	.cout());
defparam \sample_state~0 .lut_mask = 16'hAAFF;
defparam \sample_state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~1 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~1_combout ),
	.cout());
defparam \Equal6~1 .lut_mask = 16'hFFBF;
defparam \Equal6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~2 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~2_combout ),
	.cout());
defparam \Equal6~2 .lut_mask = 16'hFFDF;
defparam \Equal6~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~3 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~3_combout ),
	.cout());
defparam \Equal6~3 .lut_mask = 16'hFFEF;
defparam \Equal6~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~4 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~4_combout ),
	.cout());
defparam \Equal6~4 .lut_mask = 16'hFF7F;
defparam \Equal6~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~5 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~5_combout ),
	.cout());
defparam \Equal6~5 .lut_mask = 16'hFFFB;
defparam \Equal6~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~6 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~6_combout ),
	.cout());
defparam \Equal6~6 .lut_mask = 16'hFFFD;
defparam \Equal6~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(\ena_sample~q ),
	.datab(\Equal6~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'hEEEE;
defparam \always5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~7 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~7_combout ),
	.cout());
defparam \Equal6~7 .lut_mask = 16'hFFF7;
defparam \Equal6~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~8 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~8_combout ),
	.cout());
defparam \Equal6~8 .lut_mask = 16'hFDFF;
defparam \Equal6~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~9 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~9_combout ),
	.cout());
defparam \Equal6~9 .lut_mask = 16'hFBFF;
defparam \Equal6~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~10 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~10_combout ),
	.cout());
defparam \Equal6~10 .lut_mask = 16'hFEFF;
defparam \Equal6~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~11 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~11_combout ),
	.cout());
defparam \Equal6~11 .lut_mask = 16'hF7FF;
defparam \Equal6~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~12 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~12_combout ),
	.cout());
defparam \Equal6~12 .lut_mask = 16'hDFFF;
defparam \Equal6~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~13 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~13_combout ),
	.cout());
defparam \Equal6~13 .lut_mask = 16'hBFFF;
defparam \Equal6~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~14 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~14_combout ),
	.cout());
defparam \Equal6~14 .lut_mask = 16'hEFFF;
defparam \Equal6~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~15 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\int_channel_cnt_inst|count[2]~q ),
	.datac(\int_channel_cnt_inst|count[0]~q ),
	.datad(\int_channel_cnt_inst|count[1]~q ),
	.cin(gnd),
	.combout(\Equal6~15_combout ),
	.cout());
defparam \Equal6~15 .lut_mask = 16'h7FFF;
defparam \Equal6~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[54]~96 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[4]~6_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[46]~103_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[54]~96_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[54]~96 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[54]~96 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[53]~97 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[3]~4_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[45]~104_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[53]~97_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[53]~97 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[53]~97 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[52]~98 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[2]~2_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[44]~105_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[52]~98_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[52]~98 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[52]~98 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[61]~99 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[4]~6_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[53]~97_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[61]~99_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[61]~99 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[61]~99 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[60]~100 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[3]~4_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[52]~98_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[60]~100_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[60]~100 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[60]~100 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[59]~101 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[2]~2_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datac(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[51]~106_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[59]~101_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[59]~101 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[59]~101 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[47]~102 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[4]~6_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[8]~q ),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[47]~102_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[47]~102 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[47]~102 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[46]~103 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[3]~4_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[7]~q ),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[46]~103_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[46]~103 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[46]~103 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[45]~104 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[2]~2_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[45]~104_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[45]~104 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[45]~104 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[44]~105 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[1]~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_5_result_int[6]~10_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[44]~105_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[44]~105 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[44]~105 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[51]~106 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[1]~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_6_result_int[7]~12_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[51]~106_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[51]~106 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[51]~106 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[58]~107 (
	.dataa(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[1]~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|add_sub_7_result_int[7]~12_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datad(\Mod0|auto_generated|divider|divider|add_sub_8_result_int[7]~12_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[58]~107_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[58]~107 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[58]~107 .sum_lutc_input = "datac";

dffeas \state[0] (
	.clk(clk),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(state_0),
	.prn(vcc));
defparam \state[0] .is_wysiwyg = "true";
defparam \state[0] .power_up = "low";

dffeas \channel_out_int[0] (
	.clk(clk),
	.d(\channel_out_int~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[3]~1_combout ),
	.q(channel_out_int_0),
	.prn(vcc));
defparam \channel_out_int[0] .is_wysiwyg = "true";
defparam \channel_out_int[0] .power_up = "low";

dffeas \channel_out_int[1] (
	.clk(clk),
	.d(\channel_out_int~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[3]~1_combout ),
	.q(channel_out_int_1),
	.prn(vcc));
defparam \channel_out_int[1] .is_wysiwyg = "true";
defparam \channel_out_int[1] .power_up = "low";

dffeas \channel_out_int[2] (
	.clk(clk),
	.d(\channel_out_int~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[3]~1_combout ),
	.q(channel_out_int_2),
	.prn(vcc));
defparam \channel_out_int[2] .is_wysiwyg = "true";
defparam \channel_out_int[2] .power_up = "low";

dffeas \channel_out_int[3] (
	.clk(clk),
	.d(\channel_out_int~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[3]~1_combout ),
	.q(channel_out_int_3),
	.prn(vcc));
defparam \channel_out_int[3] .is_wysiwyg = "true";
defparam \channel_out_int[3] .power_up = "low";

cycloneive_lcell_comb \latency_cnt[2]~0 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(\state~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\latency_cnt[2]~0_combout ),
	.cout());
defparam \latency_cnt[2]~0 .lut_mask = 16'hFEFE;
defparam \latency_cnt[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \latency_cnt[0]~3 (
	.dataa(stall_reg),
	.datab(\latency_cnt[0]~q ),
	.datac(\state~0_combout ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\latency_cnt[0]~3_combout ),
	.cout());
defparam \latency_cnt[0]~3 .lut_mask = 16'h6FFF;
defparam \latency_cnt[0]~3 .sum_lutc_input = "datac";

dffeas \latency_cnt[0] (
	.clk(clk),
	.d(\latency_cnt[0]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\latency_cnt[0]~q ),
	.prn(vcc));
defparam \latency_cnt[0] .is_wysiwyg = "true";
defparam \latency_cnt[0] .power_up = "low";

cycloneive_lcell_comb \latency_cnt[1]~2 (
	.dataa(\latency_cnt[1]~q ),
	.datab(\latency_cnt[2]~0_combout ),
	.datac(reset_n),
	.datad(\latency_cnt[0]~q ),
	.cin(gnd),
	.combout(\latency_cnt[1]~2_combout ),
	.cout());
defparam \latency_cnt[1]~2 .lut_mask = 16'hF9F6;
defparam \latency_cnt[1]~2 .sum_lutc_input = "datac";

dffeas \latency_cnt[1] (
	.clk(clk),
	.d(\latency_cnt[1]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latency_cnt[1]~q ),
	.prn(vcc));
defparam \latency_cnt[1] .is_wysiwyg = "true";
defparam \latency_cnt[1] .power_up = "low";

cycloneive_lcell_comb \Add2~0 (
	.dataa(gnd),
	.datab(\latency_cnt[2]~q ),
	.datac(\latency_cnt[1]~q ),
	.datad(\latency_cnt[0]~q ),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'hC33C;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \latency_cnt[2]~1 (
	.dataa(\latency_cnt[2]~q ),
	.datab(reset_n),
	.datac(\Add2~0_combout ),
	.datad(\latency_cnt[2]~0_combout ),
	.cin(gnd),
	.combout(\latency_cnt[2]~1_combout ),
	.cout());
defparam \latency_cnt[2]~1 .lut_mask = 16'hFAFC;
defparam \latency_cnt[2]~1 .sum_lutc_input = "datac";

dffeas \latency_cnt[2] (
	.clk(clk),
	.d(\latency_cnt[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latency_cnt[2]~q ),
	.prn(vcc));
defparam \latency_cnt[2] .is_wysiwyg = "true";
defparam \latency_cnt[2] .power_up = "low";

cycloneive_lcell_comb \state~0 (
	.dataa(\latency_cnt[2]~q ),
	.datab(gnd),
	.datac(\latency_cnt[1]~q ),
	.datad(\latency_cnt[0]~q ),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hAFFF;
defparam \state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state~1 (
	.dataa(state_0),
	.datab(\state~0_combout ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'hEEFF;
defparam \state~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \channel_out_int~0 (
	.dataa(channel_out_int_0),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\channel_out_int~0_combout ),
	.cout());
defparam \channel_out_int~0 .lut_mask = 16'hFF55;
defparam \channel_out_int~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \channel_out_int[3]~1 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(dout_valid),
	.datad(state_0),
	.cin(gnd),
	.combout(\channel_out_int[3]~1_combout ),
	.cout());
defparam \channel_out_int[3]~1 .lut_mask = 16'hFFF7;
defparam \channel_out_int[3]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \channel_out_int[3]~2 (
	.dataa(channel_out_int_0),
	.datab(channel_out_int_1),
	.datac(channel_out_int_2),
	.datad(channel_out_int_3),
	.cin(gnd),
	.combout(\channel_out_int[3]~2_combout ),
	.cout());
defparam \channel_out_int[3]~2 .lut_mask = 16'h7FFF;
defparam \channel_out_int[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \channel_out_int~3 (
	.dataa(reset_n),
	.datab(\channel_out_int[3]~2_combout ),
	.datac(channel_out_int_0),
	.datad(channel_out_int_1),
	.cin(gnd),
	.combout(\channel_out_int~3_combout ),
	.cout());
defparam \channel_out_int~3 .lut_mask = 16'hEFFE;
defparam \channel_out_int~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~0 (
	.dataa(channel_out_int_0),
	.datab(channel_out_int_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'hEEEE;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \channel_out_int~4 (
	.dataa(reset_n),
	.datab(\channel_out_int[3]~2_combout ),
	.datac(channel_out_int_2),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\channel_out_int~4_combout ),
	.cout());
defparam \channel_out_int~4 .lut_mask = 16'hEFFE;
defparam \channel_out_int~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \channel_out_int~5 (
	.dataa(reset_n),
	.datab(channel_out_int_3),
	.datac(channel_out_int_2),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\channel_out_int~5_combout ),
	.cout());
defparam \channel_out_int~5 .lut_mask = 16'hEBBE;
defparam \channel_out_int~5 .sum_lutc_input = "datac";

endmodule

module CIC_auk_dspip_channel_buffer (
	q,
	fifo_rdreq_0,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_0;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_1 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_0(fifo_rdreq_0),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_1 (
	q,
	fifo_rdreq_0,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_0;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_0(fifo_rdreq_0),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51 (
	q,
	fifo_rdreq_0,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_0;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_0(fifo_rdreq_0),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu (
	q,
	fifo_rdreq_0,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_0;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_0),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_0),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_0),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_1 (
	q,
	fifo_rdreq_10,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_10;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_2 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_10(fifo_rdreq_10),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_2 (
	q,
	fifo_rdreq_10,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_10;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_1 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_10(fifo_rdreq_10),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_1 (
	q,
	fifo_rdreq_10,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_10;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_1 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_10(fifo_rdreq_10),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_1 (
	q,
	fifo_rdreq_10,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_10;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_1 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_1 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_1 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_1 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_10),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_10),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_10),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[10].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_1 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_1 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_1 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_2 (
	q,
	fifo_rdreq_11,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_11;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_3 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_11(fifo_rdreq_11),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_3 (
	q,
	fifo_rdreq_11,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_11;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_2 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_11(fifo_rdreq_11),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_2 (
	q,
	fifo_rdreq_11,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_11;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_2 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_11(fifo_rdreq_11),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_2 (
	q,
	fifo_rdreq_11,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_11;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_2 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_2 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_2 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_2 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_11),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_11),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_11),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_2 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[11].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_2 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_2 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_2 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_3 (
	q,
	fifo_rdreq_12,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_12;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_12(fifo_rdreq_12),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4 (
	q,
	fifo_rdreq_12,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_12;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_3 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_12(fifo_rdreq_12),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_3 (
	q,
	fifo_rdreq_12,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_12;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_3 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_12(fifo_rdreq_12),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_3 (
	q,
	fifo_rdreq_12,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_12;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_3 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_3 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_3 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_3 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_12),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_12),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_12),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_3 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[12].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_3 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_3 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_3 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_4 (
	q,
	fifo_rdreq_13,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_13;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_5 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_13(fifo_rdreq_13),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_5 (
	q,
	fifo_rdreq_13,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_13;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_4 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_13(fifo_rdreq_13),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_4 (
	q,
	fifo_rdreq_13,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_13;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_4 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_13(fifo_rdreq_13),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_4 (
	q,
	fifo_rdreq_13,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_13;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_4 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_4 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_4 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_4 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_13),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_13),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_13),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_4 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[13].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_4 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_4 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_4 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_5 (
	q,
	fifo_rdreq_14,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_14;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_6 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_14(fifo_rdreq_14),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_6 (
	q,
	fifo_rdreq_14,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_14;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_5 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_14(fifo_rdreq_14),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_5 (
	q,
	fifo_rdreq_14,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_14;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_5 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_14(fifo_rdreq_14),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_5 (
	q,
	fifo_rdreq_14,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_14;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_5 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_5 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_5 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_5 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_14),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_14),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_14),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_5 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[14].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_5 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_5 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_5 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_6 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_15,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_15;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_7 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_15(fifo_rdreq_15),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_7 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_15,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_15;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_6 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_15(fifo_rdreq_15),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_6 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_15,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_15;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_6 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_15(fifo_rdreq_15),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_6 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_15,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_15;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_6 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_6 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_6 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_6 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_15),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(fifo_rdreq_15),
	.datac(\empty_dff~q ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_15),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_6 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[15].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_6 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_6 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_6 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_7 (
	q,
	count_3,
	count_4,
	count_2,
	count_5,
	count_6,
	count_7,
	count_8,
	count_9,
	count_1,
	fifo_rdreq_1,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	count_3;
input 	count_4;
input 	count_2;
input 	count_5;
input 	count_6;
input 	count_7;
input 	count_8;
input 	count_9;
input 	count_1;
input 	fifo_rdreq_1;
input 	[21:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_8 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.count_3(count_3),
	.count_4(count_4),
	.count_2(count_2),
	.count_5(count_5),
	.count_6(count_6),
	.count_7(count_7),
	.count_8(count_8),
	.count_9(count_9),
	.count_1(count_1),
	.fifo_rdreq_1(fifo_rdreq_1),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.ena_sample(ena_sample),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_8 (
	q,
	count_3,
	count_4,
	count_2,
	count_5,
	count_6,
	count_7,
	count_8,
	count_9,
	count_1,
	fifo_rdreq_1,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	count_3;
input 	count_4;
input 	count_2;
input 	count_5;
input 	count_6;
input 	count_7;
input 	count_8;
input 	count_9;
input 	count_1;
input 	fifo_rdreq_1;
input 	[257:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_7 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.count_3(count_3),
	.count_4(count_4),
	.count_2(count_2),
	.count_5(count_5),
	.count_6(count_6),
	.count_7(count_7),
	.count_8(count_8),
	.count_9(count_9),
	.count_1(count_1),
	.fifo_rdreq_1(fifo_rdreq_1),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.ena_sample(ena_sample),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_7 (
	q,
	count_3,
	count_4,
	count_2,
	count_5,
	count_6,
	count_7,
	count_8,
	count_9,
	count_1,
	fifo_rdreq_1,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	count_3;
input 	count_4;
input 	count_2;
input 	count_5;
input 	count_6;
input 	count_7;
input 	count_8;
input 	count_9;
input 	count_1;
input 	fifo_rdreq_1;
input 	[21:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_7 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.count_3(count_3),
	.count_4(count_4),
	.count_2(count_2),
	.count_5(count_5),
	.count_6(count_6),
	.count_7(count_7),
	.count_8(count_8),
	.count_9(count_9),
	.count_1(count_1),
	.fifo_rdreq_1(fifo_rdreq_1),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.ena_sample(ena_sample),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_7 (
	q,
	count_3,
	count_4,
	count_2,
	count_5,
	count_6,
	count_7,
	count_8,
	count_9,
	count_1,
	fifo_rdreq_1,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	count_3;
input 	count_4;
input 	count_2;
input 	count_5;
input 	count_6;
input 	count_7;
input 	count_8;
input 	count_9;
input 	count_1;
input 	fifo_rdreq_1;
input 	[21:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~3_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;
wire \valid_wreq~0_combout ;
wire \valid_wreq~1_combout ;


CIC_cntr_u9b_7 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_7 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~3_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_7 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_7 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~3_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~3 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~3_combout ),
	.cout());
defparam \valid_wreq~3 .lut_mask = 16'hAAFF;
defparam \valid_wreq~3 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_1),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~3_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~3_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_1),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~3_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~3_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_1),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_wreq~2 (
	.dataa(ena_sample),
	.datab(\valid_wreq~0_combout ),
	.datac(\valid_wreq~1_combout ),
	.datad(count_1),
	.cin(gnd),
	.combout(valid_wreq),
	.cout());
defparam \valid_wreq~2 .lut_mask = 16'hFEFF;
defparam \valid_wreq~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(count_3),
	.datab(count_4),
	.datac(count_2),
	.datad(count_5),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'h7FFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_wreq~1 (
	.dataa(count_6),
	.datab(count_7),
	.datac(count_8),
	.datad(count_9),
	.cin(gnd),
	.combout(\valid_wreq~1_combout ),
	.cout());
defparam \valid_wreq~1 .lut_mask = 16'h7FFF;
defparam \valid_wreq~1 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_7 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_7 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_7 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_7 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_8 (
	q,
	fifo_rdreq_2,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_2;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_9 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_2(fifo_rdreq_2),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_9 (
	q,
	fifo_rdreq_2,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_2;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_8 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_2(fifo_rdreq_2),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_8 (
	q,
	fifo_rdreq_2,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_2;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_8 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_2(fifo_rdreq_2),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_8 (
	q,
	fifo_rdreq_2,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_2;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;
wire \usedw_will_be_1~3_combout ;


CIC_cntr_u9b_8 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_8 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_8 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_8 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_2),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_will_be_1~1_combout ),
	.datab(\valid_wreq~0_combout ),
	.datac(\valid_rreq~0_combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hEFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_2),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEEE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_8 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_8 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_8 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_8 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_9 (
	q,
	fifo_rdreq_3,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_3;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_10 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_3(fifo_rdreq_3),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_10 (
	q,
	fifo_rdreq_3,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_3;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_9 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_3(fifo_rdreq_3),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_9 (
	q,
	fifo_rdreq_3,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_3;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_9 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_3(fifo_rdreq_3),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_9 (
	q,
	fifo_rdreq_3,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_3;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_9 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_9 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_9 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_9 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_3),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_3),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_3),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_9 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_9 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_9 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_9 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_10 (
	q,
	fifo_rdreq_4,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_4;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_11 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_4(fifo_rdreq_4),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_11 (
	q,
	fifo_rdreq_4,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_4;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_10 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_4(fifo_rdreq_4),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_10 (
	q,
	fifo_rdreq_4,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_4;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_10 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_4(fifo_rdreq_4),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_10 (
	q,
	fifo_rdreq_4,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_4;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_10 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_10 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_10 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_10 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_4),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_4),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_4),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_10 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_10 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_10 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_10 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_11 (
	q,
	fifo_rdreq_5,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_5;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_12 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_5(fifo_rdreq_5),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_12 (
	q,
	fifo_rdreq_5,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_5;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_11 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_5(fifo_rdreq_5),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_11 (
	q,
	fifo_rdreq_5,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_5;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_11 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_5(fifo_rdreq_5),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_11 (
	q,
	fifo_rdreq_5,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_5;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_11 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_11 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_11 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_11 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_5),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_5),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_5),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_11 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_11 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_11 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_11 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_12 (
	q,
	fifo_rdreq_6,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_6;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_13 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_6(fifo_rdreq_6),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_13 (
	q,
	fifo_rdreq_6,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_6;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_12 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_6(fifo_rdreq_6),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_12 (
	q,
	fifo_rdreq_6,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_6;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_12 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_6(fifo_rdreq_6),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_12 (
	q,
	fifo_rdreq_6,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_6;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_12 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_12 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_12 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_12 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_6),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_6),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_6),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_12 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_12 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_12 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_12 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_13 (
	q,
	fifo_rdreq_7,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_7;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_14 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_7(fifo_rdreq_7),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_14 (
	q,
	fifo_rdreq_7,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_7;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_13 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_7(fifo_rdreq_7),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_13 (
	q,
	fifo_rdreq_7,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_7;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_13 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_7(fifo_rdreq_7),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_13 (
	q,
	fifo_rdreq_7,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_7;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_13 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_13 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_13 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_13 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_7),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_7),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_7),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_13 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_13 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_13 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_13 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_14 (
	q,
	fifo_rdreq_8,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_8;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_15 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_8(fifo_rdreq_8),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_15 (
	q,
	fifo_rdreq_8,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_8;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_14 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_8(fifo_rdreq_8),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_14 (
	q,
	fifo_rdreq_8,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_8;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_14 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_8(fifo_rdreq_8),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_14 (
	q,
	fifo_rdreq_8,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_8;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_14 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_14 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_14 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_14 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_8),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_8),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_8),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_14 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_14 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_14 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_14 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_channel_buffer_15 (
	q,
	fifo_rdreq_9,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_9;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_16 buffer_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,
q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_9(fifo_rdreq_9),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],
data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_16 (
	q,
	fifo_rdreq_9,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	fifo_rdreq_9;
input 	[257:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_4o51_15 auto_generated(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_9(fifo_rdreq_9),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_scfifo_4o51_15 (
	q,
	fifo_rdreq_9,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_9;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_a_dpfifo_flu_15 dpfifo(
	.q({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_unconnected_wire_4,q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.fifo_rdreq_9(fifo_rdreq_9),
	.data({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module CIC_a_dpfifo_flu_15 (
	q,
	fifo_rdreq_9,
	data,
	stall_reg,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q;
input 	fifo_rdreq_9;
input 	[21:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \usedw_counter|counter_reg_bit[4]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;


CIC_cntr_u9b_15 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_15 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_15 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_9ah1_15 FIFOram(
	.q_b({q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.data_a({data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],gnd,gnd,gnd,gnd,gnd}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_9),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAAFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(\usedw_counter|counter_reg_bit[2]~q ),
	.datab(\_~0_combout ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFFFE;
defparam \_~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~2 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~1_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hFEFF;
defparam \_~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(\_~0_combout ),
	.datab(\usedw_counter|counter_reg_bit[2]~q ),
	.datac(\usedw_counter|counter_reg_bit[4]~q ),
	.datad(\usedw_counter|counter_reg_bit[3]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(\empty_dff~q ),
	.datac(fifo_rdreq_9),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(fifo_rdreq_9),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_9ah1_15 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[21:0] q_b;
input 	[21:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 22;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 22;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 22;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 22;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 22;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 22;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 22;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 22;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 22;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 22;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 22;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 22;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 22;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 22;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 22;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 22;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 22;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 22;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 22;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 22;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 22;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 22;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 22;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 22;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 22;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 22;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 22;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 22;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 22;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 22;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 22;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 22;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[9].fifo_regulator|scfifo:buffer_FIFO|scfifo_4o51:auto_generated|a_dpfifo_flu:dpfifo|altsyncram_9ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 22;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 22;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_15 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_15 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_15 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_differentiator (
	dout_1,
	dout_2,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	stall_reg,
	dout_valid1,
	ena_diff_s_1,
	register_fifofifo_data013,
	Mux15,
	Mux16,
	Mux14,
	Mux13,
	Mux12,
	Mux11,
	Mux10,
	Mux9,
	Mux8,
	Mux7,
	Mux6,
	Mux5,
	Mux4,
	Mux3,
	Mux2,
	Mux1,
	Mux0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_1;
output 	dout_2;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
input 	stall_reg;
output 	dout_valid1;
input 	ena_diff_s_1;
input 	register_fifofifo_data013;
input 	Mux15;
input 	Mux16;
input 	Mux14;
input 	Mux13;
input 	Mux12;
input 	Mux11;
input 	Mux10;
input 	Mux9;
input 	Mux8;
input 	Mux7;
input 	Mux6;
input 	Mux5;
input 	Mux4;
input 	Mux3;
input 	Mux2;
input 	Mux1;
input 	Mux0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[15][1]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][0]~q ;
wire \glogic:u0|register_fifo:fifo_data[14][14]~0_combout ;
wire \glogic:u0|register_fifo:fifo_data[15][2]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][3]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][4]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][5]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][6]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][7]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][8]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][9]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][10]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][11]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][12]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][13]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][14]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][15]~q ;
wire \glogic:u0|register_fifo:fifo_data[15][16]~q ;
wire \dout[1]~17_cout ;
wire \dout[1]~18_combout ;
wire \dout[1]~19 ;
wire \dout[2]~20_combout ;
wire \dout[2]~21 ;
wire \dout[3]~22_combout ;
wire \dout[3]~23 ;
wire \dout[4]~24_combout ;
wire \dout[4]~25 ;
wire \dout[5]~26_combout ;
wire \dout[5]~27 ;
wire \dout[6]~28_combout ;
wire \dout[6]~29 ;
wire \dout[7]~30_combout ;
wire \dout[7]~31 ;
wire \dout[8]~32_combout ;
wire \dout[8]~33 ;
wire \dout[9]~34_combout ;
wire \dout[9]~35 ;
wire \dout[10]~36_combout ;
wire \dout[10]~37 ;
wire \dout[11]~38_combout ;
wire \dout[11]~39 ;
wire \dout[12]~40_combout ;
wire \dout[12]~41 ;
wire \dout[13]~42_combout ;
wire \dout[13]~43 ;
wire \dout[14]~44_combout ;
wire \dout[14]~45 ;
wire \dout[15]~46_combout ;
wire \dout[15]~47 ;
wire \dout[16]~48_combout ;
wire \dout_valid~0_combout ;


CIC_auk_dspip_delay \glogic:u0 (
	.stall_reg(stall_reg),
	.ena_diff_s_1(ena_diff_s_1),
	.Mux15(Mux15),
	.register_fifofifo_data151(\glogic:u0|register_fifo:fifo_data[15][1]~q ),
	.Mux16(Mux16),
	.register_fifofifo_data150(\glogic:u0|register_fifo:fifo_data[15][0]~q ),
	.register_fifofifo_data1414(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.Mux14(Mux14),
	.register_fifofifo_data152(\glogic:u0|register_fifo:fifo_data[15][2]~q ),
	.Mux13(Mux13),
	.register_fifofifo_data153(\glogic:u0|register_fifo:fifo_data[15][3]~q ),
	.Mux12(Mux12),
	.register_fifofifo_data154(\glogic:u0|register_fifo:fifo_data[15][4]~q ),
	.Mux11(Mux11),
	.register_fifofifo_data155(\glogic:u0|register_fifo:fifo_data[15][5]~q ),
	.Mux10(Mux10),
	.register_fifofifo_data156(\glogic:u0|register_fifo:fifo_data[15][6]~q ),
	.Mux9(Mux9),
	.register_fifofifo_data157(\glogic:u0|register_fifo:fifo_data[15][7]~q ),
	.Mux8(Mux8),
	.register_fifofifo_data158(\glogic:u0|register_fifo:fifo_data[15][8]~q ),
	.Mux7(Mux7),
	.register_fifofifo_data159(\glogic:u0|register_fifo:fifo_data[15][9]~q ),
	.Mux6(Mux6),
	.register_fifofifo_data1510(\glogic:u0|register_fifo:fifo_data[15][10]~q ),
	.Mux5(Mux5),
	.register_fifofifo_data1511(\glogic:u0|register_fifo:fifo_data[15][11]~q ),
	.Mux4(Mux4),
	.register_fifofifo_data1512(\glogic:u0|register_fifo:fifo_data[15][12]~q ),
	.Mux3(Mux3),
	.register_fifofifo_data1513(\glogic:u0|register_fifo:fifo_data[15][13]~q ),
	.Mux2(Mux2),
	.register_fifofifo_data1514(\glogic:u0|register_fifo:fifo_data[15][14]~q ),
	.Mux1(Mux1),
	.register_fifofifo_data1515(\glogic:u0|register_fifo:fifo_data[15][15]~q ),
	.Mux0(Mux0),
	.register_fifofifo_data1516(\glogic:u0|register_fifo:fifo_data[15][16]~q ),
	.clk(clk),
	.reset_n(reset_n));

dffeas \dout[1] (
	.clk(clk),
	.d(\dout[1]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\dout[2]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\dout[3]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\dout[4]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\dout[5]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\dout[6]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\dout[7]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\dout[8]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\dout[9]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\dout[10]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\dout[11]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\dout[12]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\dout[13]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\dout[14]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\dout[15]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\dout[16]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\glogic:u0|register_fifo:fifo_data[14][14]~0_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas dout_valid(
	.clk(clk),
	.d(\dout_valid~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data013),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

cycloneive_lcell_comb \dout[1]~17 (
	.dataa(Mux16),
	.datab(\glogic:u0|register_fifo:fifo_data[15][0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\dout[1]~17_cout ));
defparam \dout[1]~17 .lut_mask = 16'h00BB;
defparam \dout[1]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dout[1]~18 (
	.dataa(Mux15),
	.datab(\glogic:u0|register_fifo:fifo_data[15][1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[1]~17_cout ),
	.combout(\dout[1]~18_combout ),
	.cout(\dout[1]~19 ));
defparam \dout[1]~18 .lut_mask = 16'h96DF;
defparam \dout[1]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[2]~20 (
	.dataa(Mux14),
	.datab(\glogic:u0|register_fifo:fifo_data[15][2]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[1]~19 ),
	.combout(\dout[2]~20_combout ),
	.cout(\dout[2]~21 ));
defparam \dout[2]~20 .lut_mask = 16'h96BF;
defparam \dout[2]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[3]~22 (
	.dataa(Mux13),
	.datab(\glogic:u0|register_fifo:fifo_data[15][3]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[2]~21 ),
	.combout(\dout[3]~22_combout ),
	.cout(\dout[3]~23 ));
defparam \dout[3]~22 .lut_mask = 16'h96DF;
defparam \dout[3]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[4]~24 (
	.dataa(Mux12),
	.datab(\glogic:u0|register_fifo:fifo_data[15][4]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[3]~23 ),
	.combout(\dout[4]~24_combout ),
	.cout(\dout[4]~25 ));
defparam \dout[4]~24 .lut_mask = 16'h96BF;
defparam \dout[4]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[5]~26 (
	.dataa(Mux11),
	.datab(\glogic:u0|register_fifo:fifo_data[15][5]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[4]~25 ),
	.combout(\dout[5]~26_combout ),
	.cout(\dout[5]~27 ));
defparam \dout[5]~26 .lut_mask = 16'h96DF;
defparam \dout[5]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[6]~28 (
	.dataa(Mux10),
	.datab(\glogic:u0|register_fifo:fifo_data[15][6]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[5]~27 ),
	.combout(\dout[6]~28_combout ),
	.cout(\dout[6]~29 ));
defparam \dout[6]~28 .lut_mask = 16'h96BF;
defparam \dout[6]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[7]~30 (
	.dataa(Mux9),
	.datab(\glogic:u0|register_fifo:fifo_data[15][7]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[6]~29 ),
	.combout(\dout[7]~30_combout ),
	.cout(\dout[7]~31 ));
defparam \dout[7]~30 .lut_mask = 16'h96DF;
defparam \dout[7]~30 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[8]~32 (
	.dataa(Mux8),
	.datab(\glogic:u0|register_fifo:fifo_data[15][8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[7]~31 ),
	.combout(\dout[8]~32_combout ),
	.cout(\dout[8]~33 ));
defparam \dout[8]~32 .lut_mask = 16'h96BF;
defparam \dout[8]~32 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[9]~34 (
	.dataa(Mux7),
	.datab(\glogic:u0|register_fifo:fifo_data[15][9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[8]~33 ),
	.combout(\dout[9]~34_combout ),
	.cout(\dout[9]~35 ));
defparam \dout[9]~34 .lut_mask = 16'h96DF;
defparam \dout[9]~34 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[10]~36 (
	.dataa(Mux6),
	.datab(\glogic:u0|register_fifo:fifo_data[15][10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[9]~35 ),
	.combout(\dout[10]~36_combout ),
	.cout(\dout[10]~37 ));
defparam \dout[10]~36 .lut_mask = 16'h96BF;
defparam \dout[10]~36 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[11]~38 (
	.dataa(Mux5),
	.datab(\glogic:u0|register_fifo:fifo_data[15][11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[10]~37 ),
	.combout(\dout[11]~38_combout ),
	.cout(\dout[11]~39 ));
defparam \dout[11]~38 .lut_mask = 16'h96DF;
defparam \dout[11]~38 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[12]~40 (
	.dataa(Mux4),
	.datab(\glogic:u0|register_fifo:fifo_data[15][12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[11]~39 ),
	.combout(\dout[12]~40_combout ),
	.cout(\dout[12]~41 ));
defparam \dout[12]~40 .lut_mask = 16'h96BF;
defparam \dout[12]~40 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[13]~42 (
	.dataa(Mux3),
	.datab(\glogic:u0|register_fifo:fifo_data[15][13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[12]~41 ),
	.combout(\dout[13]~42_combout ),
	.cout(\dout[13]~43 ));
defparam \dout[13]~42 .lut_mask = 16'h96DF;
defparam \dout[13]~42 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[14]~44 (
	.dataa(Mux2),
	.datab(\glogic:u0|register_fifo:fifo_data[15][14]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[13]~43 ),
	.combout(\dout[14]~44_combout ),
	.cout(\dout[14]~45 ));
defparam \dout[14]~44 .lut_mask = 16'h96BF;
defparam \dout[14]~44 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[15]~46 (
	.dataa(Mux1),
	.datab(\glogic:u0|register_fifo:fifo_data[15][15]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[14]~45 ),
	.combout(\dout[15]~46_combout ),
	.cout(\dout[15]~47 ));
defparam \dout[15]~46 .lut_mask = 16'h96DF;
defparam \dout[15]~46 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout[16]~48 (
	.dataa(Mux0),
	.datab(\glogic:u0|register_fifo:fifo_data[15][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dout[15]~47 ),
	.combout(\dout[16]~48_combout ),
	.cout());
defparam \dout[16]~48 .lut_mask = 16'h9696;
defparam \dout[16]~48 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dout_valid~0 (
	.dataa(reset_n),
	.datab(ena_diff_s_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dout_valid~0_combout ),
	.cout());
defparam \dout_valid~0 .lut_mask = 16'hEEEE;
defparam \dout_valid~0 .sum_lutc_input = "datac";

endmodule

module CIC_auk_dspip_delay (
	stall_reg,
	ena_diff_s_1,
	Mux15,
	register_fifofifo_data151,
	Mux16,
	register_fifofifo_data150,
	register_fifofifo_data1414,
	Mux14,
	register_fifofifo_data152,
	Mux13,
	register_fifofifo_data153,
	Mux12,
	register_fifofifo_data154,
	Mux11,
	register_fifofifo_data155,
	Mux10,
	register_fifofifo_data156,
	Mux9,
	register_fifofifo_data157,
	Mux8,
	register_fifofifo_data158,
	Mux7,
	register_fifofifo_data159,
	Mux6,
	register_fifofifo_data1510,
	Mux5,
	register_fifofifo_data1511,
	Mux4,
	register_fifofifo_data1512,
	Mux3,
	register_fifofifo_data1513,
	Mux2,
	register_fifofifo_data1514,
	Mux1,
	register_fifofifo_data1515,
	Mux0,
	register_fifofifo_data1516,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	stall_reg;
input 	ena_diff_s_1;
input 	Mux15;
output 	register_fifofifo_data151;
input 	Mux16;
output 	register_fifofifo_data150;
output 	register_fifofifo_data1414;
input 	Mux14;
output 	register_fifofifo_data152;
input 	Mux13;
output 	register_fifofifo_data153;
input 	Mux12;
output 	register_fifofifo_data154;
input 	Mux11;
output 	register_fifofifo_data155;
input 	Mux10;
output 	register_fifofifo_data156;
input 	Mux9;
output 	register_fifofifo_data157;
input 	Mux8;
output 	register_fifofifo_data158;
input 	Mux7;
output 	register_fifofifo_data159;
input 	Mux6;
output 	register_fifofifo_data1510;
input 	Mux5;
output 	register_fifofifo_data1511;
input 	Mux4;
output 	register_fifofifo_data1512;
input 	Mux3;
output 	register_fifofifo_data1513;
input 	Mux2;
output 	register_fifofifo_data1514;
input 	Mux1;
output 	register_fifofifo_data1515;
input 	Mux0;
output 	register_fifofifo_data1516;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fifo_data~255_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \fifo_data~238_combout ;
wire \register_fifo:fifo_data[1][1]~q ;
wire \fifo_data~221_combout ;
wire \register_fifo:fifo_data[2][1]~q ;
wire \fifo_data~204_combout ;
wire \register_fifo:fifo_data[3][1]~q ;
wire \fifo_data~187_combout ;
wire \register_fifo:fifo_data[4][1]~q ;
wire \fifo_data~170_combout ;
wire \register_fifo:fifo_data[5][1]~q ;
wire \fifo_data~153_combout ;
wire \register_fifo:fifo_data[6][1]~q ;
wire \fifo_data~136_combout ;
wire \register_fifo:fifo_data[7][1]~q ;
wire \fifo_data~119_combout ;
wire \register_fifo:fifo_data[8][1]~q ;
wire \fifo_data~102_combout ;
wire \register_fifo:fifo_data[9][1]~q ;
wire \fifo_data~85_combout ;
wire \register_fifo:fifo_data[10][1]~q ;
wire \fifo_data~68_combout ;
wire \register_fifo:fifo_data[11][1]~q ;
wire \fifo_data~51_combout ;
wire \register_fifo:fifo_data[12][1]~q ;
wire \fifo_data~34_combout ;
wire \register_fifo:fifo_data[13][1]~q ;
wire \fifo_data~17_combout ;
wire \register_fifo:fifo_data[14][1]~q ;
wire \fifo_data~0_combout ;
wire \fifo_data~256_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \fifo_data~239_combout ;
wire \register_fifo:fifo_data[1][0]~q ;
wire \fifo_data~222_combout ;
wire \register_fifo:fifo_data[2][0]~q ;
wire \fifo_data~205_combout ;
wire \register_fifo:fifo_data[3][0]~q ;
wire \fifo_data~188_combout ;
wire \register_fifo:fifo_data[4][0]~q ;
wire \fifo_data~171_combout ;
wire \register_fifo:fifo_data[5][0]~q ;
wire \fifo_data~154_combout ;
wire \register_fifo:fifo_data[6][0]~q ;
wire \fifo_data~137_combout ;
wire \register_fifo:fifo_data[7][0]~q ;
wire \fifo_data~120_combout ;
wire \register_fifo:fifo_data[8][0]~q ;
wire \fifo_data~103_combout ;
wire \register_fifo:fifo_data[9][0]~q ;
wire \fifo_data~86_combout ;
wire \register_fifo:fifo_data[10][0]~q ;
wire \fifo_data~69_combout ;
wire \register_fifo:fifo_data[11][0]~q ;
wire \fifo_data~52_combout ;
wire \register_fifo:fifo_data[12][0]~q ;
wire \fifo_data~35_combout ;
wire \register_fifo:fifo_data[13][0]~q ;
wire \fifo_data~18_combout ;
wire \register_fifo:fifo_data[14][0]~q ;
wire \fifo_data~1_combout ;
wire \fifo_data~257_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \fifo_data~240_combout ;
wire \register_fifo:fifo_data[1][2]~q ;
wire \fifo_data~223_combout ;
wire \register_fifo:fifo_data[2][2]~q ;
wire \fifo_data~206_combout ;
wire \register_fifo:fifo_data[3][2]~q ;
wire \fifo_data~189_combout ;
wire \register_fifo:fifo_data[4][2]~q ;
wire \fifo_data~172_combout ;
wire \register_fifo:fifo_data[5][2]~q ;
wire \fifo_data~155_combout ;
wire \register_fifo:fifo_data[6][2]~q ;
wire \fifo_data~138_combout ;
wire \register_fifo:fifo_data[7][2]~q ;
wire \fifo_data~121_combout ;
wire \register_fifo:fifo_data[8][2]~q ;
wire \fifo_data~104_combout ;
wire \register_fifo:fifo_data[9][2]~q ;
wire \fifo_data~87_combout ;
wire \register_fifo:fifo_data[10][2]~q ;
wire \fifo_data~70_combout ;
wire \register_fifo:fifo_data[11][2]~q ;
wire \fifo_data~53_combout ;
wire \register_fifo:fifo_data[12][2]~q ;
wire \fifo_data~36_combout ;
wire \register_fifo:fifo_data[13][2]~q ;
wire \fifo_data~19_combout ;
wire \register_fifo:fifo_data[14][2]~q ;
wire \fifo_data~2_combout ;
wire \fifo_data~258_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \fifo_data~241_combout ;
wire \register_fifo:fifo_data[1][3]~q ;
wire \fifo_data~224_combout ;
wire \register_fifo:fifo_data[2][3]~q ;
wire \fifo_data~207_combout ;
wire \register_fifo:fifo_data[3][3]~q ;
wire \fifo_data~190_combout ;
wire \register_fifo:fifo_data[4][3]~q ;
wire \fifo_data~173_combout ;
wire \register_fifo:fifo_data[5][3]~q ;
wire \fifo_data~156_combout ;
wire \register_fifo:fifo_data[6][3]~q ;
wire \fifo_data~139_combout ;
wire \register_fifo:fifo_data[7][3]~q ;
wire \fifo_data~122_combout ;
wire \register_fifo:fifo_data[8][3]~q ;
wire \fifo_data~105_combout ;
wire \register_fifo:fifo_data[9][3]~q ;
wire \fifo_data~88_combout ;
wire \register_fifo:fifo_data[10][3]~q ;
wire \fifo_data~71_combout ;
wire \register_fifo:fifo_data[11][3]~q ;
wire \fifo_data~54_combout ;
wire \register_fifo:fifo_data[12][3]~q ;
wire \fifo_data~37_combout ;
wire \register_fifo:fifo_data[13][3]~q ;
wire \fifo_data~20_combout ;
wire \register_fifo:fifo_data[14][3]~q ;
wire \fifo_data~3_combout ;
wire \fifo_data~259_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \fifo_data~242_combout ;
wire \register_fifo:fifo_data[1][4]~q ;
wire \fifo_data~225_combout ;
wire \register_fifo:fifo_data[2][4]~q ;
wire \fifo_data~208_combout ;
wire \register_fifo:fifo_data[3][4]~q ;
wire \fifo_data~191_combout ;
wire \register_fifo:fifo_data[4][4]~q ;
wire \fifo_data~174_combout ;
wire \register_fifo:fifo_data[5][4]~q ;
wire \fifo_data~157_combout ;
wire \register_fifo:fifo_data[6][4]~q ;
wire \fifo_data~140_combout ;
wire \register_fifo:fifo_data[7][4]~q ;
wire \fifo_data~123_combout ;
wire \register_fifo:fifo_data[8][4]~q ;
wire \fifo_data~106_combout ;
wire \register_fifo:fifo_data[9][4]~q ;
wire \fifo_data~89_combout ;
wire \register_fifo:fifo_data[10][4]~q ;
wire \fifo_data~72_combout ;
wire \register_fifo:fifo_data[11][4]~q ;
wire \fifo_data~55_combout ;
wire \register_fifo:fifo_data[12][4]~q ;
wire \fifo_data~38_combout ;
wire \register_fifo:fifo_data[13][4]~q ;
wire \fifo_data~21_combout ;
wire \register_fifo:fifo_data[14][4]~q ;
wire \fifo_data~4_combout ;
wire \fifo_data~260_combout ;
wire \register_fifo:fifo_data[0][5]~q ;
wire \fifo_data~243_combout ;
wire \register_fifo:fifo_data[1][5]~q ;
wire \fifo_data~226_combout ;
wire \register_fifo:fifo_data[2][5]~q ;
wire \fifo_data~209_combout ;
wire \register_fifo:fifo_data[3][5]~q ;
wire \fifo_data~192_combout ;
wire \register_fifo:fifo_data[4][5]~q ;
wire \fifo_data~175_combout ;
wire \register_fifo:fifo_data[5][5]~q ;
wire \fifo_data~158_combout ;
wire \register_fifo:fifo_data[6][5]~q ;
wire \fifo_data~141_combout ;
wire \register_fifo:fifo_data[7][5]~q ;
wire \fifo_data~124_combout ;
wire \register_fifo:fifo_data[8][5]~q ;
wire \fifo_data~107_combout ;
wire \register_fifo:fifo_data[9][5]~q ;
wire \fifo_data~90_combout ;
wire \register_fifo:fifo_data[10][5]~q ;
wire \fifo_data~73_combout ;
wire \register_fifo:fifo_data[11][5]~q ;
wire \fifo_data~56_combout ;
wire \register_fifo:fifo_data[12][5]~q ;
wire \fifo_data~39_combout ;
wire \register_fifo:fifo_data[13][5]~q ;
wire \fifo_data~22_combout ;
wire \register_fifo:fifo_data[14][5]~q ;
wire \fifo_data~5_combout ;
wire \fifo_data~261_combout ;
wire \register_fifo:fifo_data[0][6]~q ;
wire \fifo_data~244_combout ;
wire \register_fifo:fifo_data[1][6]~q ;
wire \fifo_data~227_combout ;
wire \register_fifo:fifo_data[2][6]~q ;
wire \fifo_data~210_combout ;
wire \register_fifo:fifo_data[3][6]~q ;
wire \fifo_data~193_combout ;
wire \register_fifo:fifo_data[4][6]~q ;
wire \fifo_data~176_combout ;
wire \register_fifo:fifo_data[5][6]~q ;
wire \fifo_data~159_combout ;
wire \register_fifo:fifo_data[6][6]~q ;
wire \fifo_data~142_combout ;
wire \register_fifo:fifo_data[7][6]~q ;
wire \fifo_data~125_combout ;
wire \register_fifo:fifo_data[8][6]~q ;
wire \fifo_data~108_combout ;
wire \register_fifo:fifo_data[9][6]~q ;
wire \fifo_data~91_combout ;
wire \register_fifo:fifo_data[10][6]~q ;
wire \fifo_data~74_combout ;
wire \register_fifo:fifo_data[11][6]~q ;
wire \fifo_data~57_combout ;
wire \register_fifo:fifo_data[12][6]~q ;
wire \fifo_data~40_combout ;
wire \register_fifo:fifo_data[13][6]~q ;
wire \fifo_data~23_combout ;
wire \register_fifo:fifo_data[14][6]~q ;
wire \fifo_data~6_combout ;
wire \fifo_data~262_combout ;
wire \register_fifo:fifo_data[0][7]~q ;
wire \fifo_data~245_combout ;
wire \register_fifo:fifo_data[1][7]~q ;
wire \fifo_data~228_combout ;
wire \register_fifo:fifo_data[2][7]~q ;
wire \fifo_data~211_combout ;
wire \register_fifo:fifo_data[3][7]~q ;
wire \fifo_data~194_combout ;
wire \register_fifo:fifo_data[4][7]~q ;
wire \fifo_data~177_combout ;
wire \register_fifo:fifo_data[5][7]~q ;
wire \fifo_data~160_combout ;
wire \register_fifo:fifo_data[6][7]~q ;
wire \fifo_data~143_combout ;
wire \register_fifo:fifo_data[7][7]~q ;
wire \fifo_data~126_combout ;
wire \register_fifo:fifo_data[8][7]~q ;
wire \fifo_data~109_combout ;
wire \register_fifo:fifo_data[9][7]~q ;
wire \fifo_data~92_combout ;
wire \register_fifo:fifo_data[10][7]~q ;
wire \fifo_data~75_combout ;
wire \register_fifo:fifo_data[11][7]~q ;
wire \fifo_data~58_combout ;
wire \register_fifo:fifo_data[12][7]~q ;
wire \fifo_data~41_combout ;
wire \register_fifo:fifo_data[13][7]~q ;
wire \fifo_data~24_combout ;
wire \register_fifo:fifo_data[14][7]~q ;
wire \fifo_data~7_combout ;
wire \fifo_data~263_combout ;
wire \register_fifo:fifo_data[0][8]~q ;
wire \fifo_data~246_combout ;
wire \register_fifo:fifo_data[1][8]~q ;
wire \fifo_data~229_combout ;
wire \register_fifo:fifo_data[2][8]~q ;
wire \fifo_data~212_combout ;
wire \register_fifo:fifo_data[3][8]~q ;
wire \fifo_data~195_combout ;
wire \register_fifo:fifo_data[4][8]~q ;
wire \fifo_data~178_combout ;
wire \register_fifo:fifo_data[5][8]~q ;
wire \fifo_data~161_combout ;
wire \register_fifo:fifo_data[6][8]~q ;
wire \fifo_data~144_combout ;
wire \register_fifo:fifo_data[7][8]~q ;
wire \fifo_data~127_combout ;
wire \register_fifo:fifo_data[8][8]~q ;
wire \fifo_data~110_combout ;
wire \register_fifo:fifo_data[9][8]~q ;
wire \fifo_data~93_combout ;
wire \register_fifo:fifo_data[10][8]~q ;
wire \fifo_data~76_combout ;
wire \register_fifo:fifo_data[11][8]~q ;
wire \fifo_data~59_combout ;
wire \register_fifo:fifo_data[12][8]~q ;
wire \fifo_data~42_combout ;
wire \register_fifo:fifo_data[13][8]~q ;
wire \fifo_data~25_combout ;
wire \register_fifo:fifo_data[14][8]~q ;
wire \fifo_data~8_combout ;
wire \fifo_data~264_combout ;
wire \register_fifo:fifo_data[0][9]~q ;
wire \fifo_data~247_combout ;
wire \register_fifo:fifo_data[1][9]~q ;
wire \fifo_data~230_combout ;
wire \register_fifo:fifo_data[2][9]~q ;
wire \fifo_data~213_combout ;
wire \register_fifo:fifo_data[3][9]~q ;
wire \fifo_data~196_combout ;
wire \register_fifo:fifo_data[4][9]~q ;
wire \fifo_data~179_combout ;
wire \register_fifo:fifo_data[5][9]~q ;
wire \fifo_data~162_combout ;
wire \register_fifo:fifo_data[6][9]~q ;
wire \fifo_data~145_combout ;
wire \register_fifo:fifo_data[7][9]~q ;
wire \fifo_data~128_combout ;
wire \register_fifo:fifo_data[8][9]~q ;
wire \fifo_data~111_combout ;
wire \register_fifo:fifo_data[9][9]~q ;
wire \fifo_data~94_combout ;
wire \register_fifo:fifo_data[10][9]~q ;
wire \fifo_data~77_combout ;
wire \register_fifo:fifo_data[11][9]~q ;
wire \fifo_data~60_combout ;
wire \register_fifo:fifo_data[12][9]~q ;
wire \fifo_data~43_combout ;
wire \register_fifo:fifo_data[13][9]~q ;
wire \fifo_data~26_combout ;
wire \register_fifo:fifo_data[14][9]~q ;
wire \fifo_data~9_combout ;
wire \fifo_data~265_combout ;
wire \register_fifo:fifo_data[0][10]~q ;
wire \fifo_data~248_combout ;
wire \register_fifo:fifo_data[1][10]~q ;
wire \fifo_data~231_combout ;
wire \register_fifo:fifo_data[2][10]~q ;
wire \fifo_data~214_combout ;
wire \register_fifo:fifo_data[3][10]~q ;
wire \fifo_data~197_combout ;
wire \register_fifo:fifo_data[4][10]~q ;
wire \fifo_data~180_combout ;
wire \register_fifo:fifo_data[5][10]~q ;
wire \fifo_data~163_combout ;
wire \register_fifo:fifo_data[6][10]~q ;
wire \fifo_data~146_combout ;
wire \register_fifo:fifo_data[7][10]~q ;
wire \fifo_data~129_combout ;
wire \register_fifo:fifo_data[8][10]~q ;
wire \fifo_data~112_combout ;
wire \register_fifo:fifo_data[9][10]~q ;
wire \fifo_data~95_combout ;
wire \register_fifo:fifo_data[10][10]~q ;
wire \fifo_data~78_combout ;
wire \register_fifo:fifo_data[11][10]~q ;
wire \fifo_data~61_combout ;
wire \register_fifo:fifo_data[12][10]~q ;
wire \fifo_data~44_combout ;
wire \register_fifo:fifo_data[13][10]~q ;
wire \fifo_data~27_combout ;
wire \register_fifo:fifo_data[14][10]~q ;
wire \fifo_data~10_combout ;
wire \fifo_data~266_combout ;
wire \register_fifo:fifo_data[0][11]~q ;
wire \fifo_data~249_combout ;
wire \register_fifo:fifo_data[1][11]~q ;
wire \fifo_data~232_combout ;
wire \register_fifo:fifo_data[2][11]~q ;
wire \fifo_data~215_combout ;
wire \register_fifo:fifo_data[3][11]~q ;
wire \fifo_data~198_combout ;
wire \register_fifo:fifo_data[4][11]~q ;
wire \fifo_data~181_combout ;
wire \register_fifo:fifo_data[5][11]~q ;
wire \fifo_data~164_combout ;
wire \register_fifo:fifo_data[6][11]~q ;
wire \fifo_data~147_combout ;
wire \register_fifo:fifo_data[7][11]~q ;
wire \fifo_data~130_combout ;
wire \register_fifo:fifo_data[8][11]~q ;
wire \fifo_data~113_combout ;
wire \register_fifo:fifo_data[9][11]~q ;
wire \fifo_data~96_combout ;
wire \register_fifo:fifo_data[10][11]~q ;
wire \fifo_data~79_combout ;
wire \register_fifo:fifo_data[11][11]~q ;
wire \fifo_data~62_combout ;
wire \register_fifo:fifo_data[12][11]~q ;
wire \fifo_data~45_combout ;
wire \register_fifo:fifo_data[13][11]~q ;
wire \fifo_data~28_combout ;
wire \register_fifo:fifo_data[14][11]~q ;
wire \fifo_data~11_combout ;
wire \fifo_data~267_combout ;
wire \register_fifo:fifo_data[0][12]~q ;
wire \fifo_data~250_combout ;
wire \register_fifo:fifo_data[1][12]~q ;
wire \fifo_data~233_combout ;
wire \register_fifo:fifo_data[2][12]~q ;
wire \fifo_data~216_combout ;
wire \register_fifo:fifo_data[3][12]~q ;
wire \fifo_data~199_combout ;
wire \register_fifo:fifo_data[4][12]~q ;
wire \fifo_data~182_combout ;
wire \register_fifo:fifo_data[5][12]~q ;
wire \fifo_data~165_combout ;
wire \register_fifo:fifo_data[6][12]~q ;
wire \fifo_data~148_combout ;
wire \register_fifo:fifo_data[7][12]~q ;
wire \fifo_data~131_combout ;
wire \register_fifo:fifo_data[8][12]~q ;
wire \fifo_data~114_combout ;
wire \register_fifo:fifo_data[9][12]~q ;
wire \fifo_data~97_combout ;
wire \register_fifo:fifo_data[10][12]~q ;
wire \fifo_data~80_combout ;
wire \register_fifo:fifo_data[11][12]~q ;
wire \fifo_data~63_combout ;
wire \register_fifo:fifo_data[12][12]~q ;
wire \fifo_data~46_combout ;
wire \register_fifo:fifo_data[13][12]~q ;
wire \fifo_data~29_combout ;
wire \register_fifo:fifo_data[14][12]~q ;
wire \fifo_data~12_combout ;
wire \fifo_data~268_combout ;
wire \register_fifo:fifo_data[0][13]~q ;
wire \fifo_data~251_combout ;
wire \register_fifo:fifo_data[1][13]~q ;
wire \fifo_data~234_combout ;
wire \register_fifo:fifo_data[2][13]~q ;
wire \fifo_data~217_combout ;
wire \register_fifo:fifo_data[3][13]~q ;
wire \fifo_data~200_combout ;
wire \register_fifo:fifo_data[4][13]~q ;
wire \fifo_data~183_combout ;
wire \register_fifo:fifo_data[5][13]~q ;
wire \fifo_data~166_combout ;
wire \register_fifo:fifo_data[6][13]~q ;
wire \fifo_data~149_combout ;
wire \register_fifo:fifo_data[7][13]~q ;
wire \fifo_data~132_combout ;
wire \register_fifo:fifo_data[8][13]~q ;
wire \fifo_data~115_combout ;
wire \register_fifo:fifo_data[9][13]~q ;
wire \fifo_data~98_combout ;
wire \register_fifo:fifo_data[10][13]~q ;
wire \fifo_data~81_combout ;
wire \register_fifo:fifo_data[11][13]~q ;
wire \fifo_data~64_combout ;
wire \register_fifo:fifo_data[12][13]~q ;
wire \fifo_data~47_combout ;
wire \register_fifo:fifo_data[13][13]~q ;
wire \fifo_data~30_combout ;
wire \register_fifo:fifo_data[14][13]~q ;
wire \fifo_data~13_combout ;
wire \fifo_data~269_combout ;
wire \register_fifo:fifo_data[0][14]~q ;
wire \fifo_data~252_combout ;
wire \register_fifo:fifo_data[1][14]~q ;
wire \fifo_data~235_combout ;
wire \register_fifo:fifo_data[2][14]~q ;
wire \fifo_data~218_combout ;
wire \register_fifo:fifo_data[3][14]~q ;
wire \fifo_data~201_combout ;
wire \register_fifo:fifo_data[4][14]~q ;
wire \fifo_data~184_combout ;
wire \register_fifo:fifo_data[5][14]~q ;
wire \fifo_data~167_combout ;
wire \register_fifo:fifo_data[6][14]~q ;
wire \fifo_data~150_combout ;
wire \register_fifo:fifo_data[7][14]~q ;
wire \fifo_data~133_combout ;
wire \register_fifo:fifo_data[8][14]~q ;
wire \fifo_data~116_combout ;
wire \register_fifo:fifo_data[9][14]~q ;
wire \fifo_data~99_combout ;
wire \register_fifo:fifo_data[10][14]~q ;
wire \fifo_data~82_combout ;
wire \register_fifo:fifo_data[11][14]~q ;
wire \fifo_data~65_combout ;
wire \register_fifo:fifo_data[12][14]~q ;
wire \fifo_data~48_combout ;
wire \register_fifo:fifo_data[13][14]~q ;
wire \fifo_data~31_combout ;
wire \register_fifo:fifo_data[14][14]~q ;
wire \fifo_data~14_combout ;
wire \fifo_data~270_combout ;
wire \register_fifo:fifo_data[0][15]~q ;
wire \fifo_data~253_combout ;
wire \register_fifo:fifo_data[1][15]~q ;
wire \fifo_data~236_combout ;
wire \register_fifo:fifo_data[2][15]~q ;
wire \fifo_data~219_combout ;
wire \register_fifo:fifo_data[3][15]~q ;
wire \fifo_data~202_combout ;
wire \register_fifo:fifo_data[4][15]~q ;
wire \fifo_data~185_combout ;
wire \register_fifo:fifo_data[5][15]~q ;
wire \fifo_data~168_combout ;
wire \register_fifo:fifo_data[6][15]~q ;
wire \fifo_data~151_combout ;
wire \register_fifo:fifo_data[7][15]~q ;
wire \fifo_data~134_combout ;
wire \register_fifo:fifo_data[8][15]~q ;
wire \fifo_data~117_combout ;
wire \register_fifo:fifo_data[9][15]~q ;
wire \fifo_data~100_combout ;
wire \register_fifo:fifo_data[10][15]~q ;
wire \fifo_data~83_combout ;
wire \register_fifo:fifo_data[11][15]~q ;
wire \fifo_data~66_combout ;
wire \register_fifo:fifo_data[12][15]~q ;
wire \fifo_data~49_combout ;
wire \register_fifo:fifo_data[13][15]~q ;
wire \fifo_data~32_combout ;
wire \register_fifo:fifo_data[14][15]~q ;
wire \fifo_data~15_combout ;
wire \fifo_data~271_combout ;
wire \register_fifo:fifo_data[0][16]~q ;
wire \fifo_data~254_combout ;
wire \register_fifo:fifo_data[1][16]~q ;
wire \fifo_data~237_combout ;
wire \register_fifo:fifo_data[2][16]~q ;
wire \fifo_data~220_combout ;
wire \register_fifo:fifo_data[3][16]~q ;
wire \fifo_data~203_combout ;
wire \register_fifo:fifo_data[4][16]~q ;
wire \fifo_data~186_combout ;
wire \register_fifo:fifo_data[5][16]~q ;
wire \fifo_data~169_combout ;
wire \register_fifo:fifo_data[6][16]~q ;
wire \fifo_data~152_combout ;
wire \register_fifo:fifo_data[7][16]~q ;
wire \fifo_data~135_combout ;
wire \register_fifo:fifo_data[8][16]~q ;
wire \fifo_data~118_combout ;
wire \register_fifo:fifo_data[9][16]~q ;
wire \fifo_data~101_combout ;
wire \register_fifo:fifo_data[10][16]~q ;
wire \fifo_data~84_combout ;
wire \register_fifo:fifo_data[11][16]~q ;
wire \fifo_data~67_combout ;
wire \register_fifo:fifo_data[12][16]~q ;
wire \fifo_data~50_combout ;
wire \register_fifo:fifo_data[13][16]~q ;
wire \fifo_data~33_combout ;
wire \register_fifo:fifo_data[14][16]~q ;
wire \fifo_data~16_combout ;


dffeas \register_fifo:fifo_data[15][1] (
	.clk(clk),
	.d(\fifo_data~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data151),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][1] .power_up = "low";

dffeas \register_fifo:fifo_data[15][0] (
	.clk(clk),
	.d(\fifo_data~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data150),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[14][14]~0 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(ena_diff_s_1),
	.cin(gnd),
	.combout(register_fifofifo_data1414),
	.cout());
defparam \register_fifo:fifo_data[14][14]~0 .lut_mask = 16'hFF77;
defparam \register_fifo:fifo_data[14][14]~0 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[15][2] (
	.clk(clk),
	.d(\fifo_data~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data152),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][2] .power_up = "low";

dffeas \register_fifo:fifo_data[15][3] (
	.clk(clk),
	.d(\fifo_data~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data153),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][3] .power_up = "low";

dffeas \register_fifo:fifo_data[15][4] (
	.clk(clk),
	.d(\fifo_data~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data154),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][4] .power_up = "low";

dffeas \register_fifo:fifo_data[15][5] (
	.clk(clk),
	.d(\fifo_data~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data155),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][5] .power_up = "low";

dffeas \register_fifo:fifo_data[15][6] (
	.clk(clk),
	.d(\fifo_data~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data156),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][6] .power_up = "low";

dffeas \register_fifo:fifo_data[15][7] (
	.clk(clk),
	.d(\fifo_data~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data157),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][7] .power_up = "low";

dffeas \register_fifo:fifo_data[15][8] (
	.clk(clk),
	.d(\fifo_data~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data158),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][8] .power_up = "low";

dffeas \register_fifo:fifo_data[15][9] (
	.clk(clk),
	.d(\fifo_data~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data159),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][9] .power_up = "low";

dffeas \register_fifo:fifo_data[15][10] (
	.clk(clk),
	.d(\fifo_data~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data1510),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][10] .power_up = "low";

dffeas \register_fifo:fifo_data[15][11] (
	.clk(clk),
	.d(\fifo_data~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data1511),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][11] .power_up = "low";

dffeas \register_fifo:fifo_data[15][12] (
	.clk(clk),
	.d(\fifo_data~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data1512),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][12] .power_up = "low";

dffeas \register_fifo:fifo_data[15][13] (
	.clk(clk),
	.d(\fifo_data~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data1513),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][13] .power_up = "low";

dffeas \register_fifo:fifo_data[15][14] (
	.clk(clk),
	.d(\fifo_data~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data1514),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][14] .power_up = "low";

dffeas \register_fifo:fifo_data[15][15] (
	.clk(clk),
	.d(\fifo_data~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data1515),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][15] .power_up = "low";

dffeas \register_fifo:fifo_data[15][16] (
	.clk(clk),
	.d(\fifo_data~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(register_fifofifo_data1516),
	.prn(vcc));
defparam \register_fifo:fifo_data[15][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[15][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~255 (
	.dataa(reset_n),
	.datab(Mux15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~255_combout ),
	.cout());
defparam \fifo_data~255 .lut_mask = 16'hEEEE;
defparam \fifo_data~255 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\fifo_data~255_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~238 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~238_combout ),
	.cout());
defparam \fifo_data~238 .lut_mask = 16'hEEEE;
defparam \fifo_data~238 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][1] (
	.clk(clk),
	.d(\fifo_data~238_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~221 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~221_combout ),
	.cout());
defparam \fifo_data~221 .lut_mask = 16'hEEEE;
defparam \fifo_data~221 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][1] (
	.clk(clk),
	.d(\fifo_data~221_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~204 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~204_combout ),
	.cout());
defparam \fifo_data~204 .lut_mask = 16'hEEEE;
defparam \fifo_data~204 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][1] (
	.clk(clk),
	.d(\fifo_data~204_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~187 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~187_combout ),
	.cout());
defparam \fifo_data~187 .lut_mask = 16'hEEEE;
defparam \fifo_data~187 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][1] (
	.clk(clk),
	.d(\fifo_data~187_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~170 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~170_combout ),
	.cout());
defparam \fifo_data~170 .lut_mask = 16'hEEEE;
defparam \fifo_data~170 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][1] (
	.clk(clk),
	.d(\fifo_data~170_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~153 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~153_combout ),
	.cout());
defparam \fifo_data~153 .lut_mask = 16'hEEEE;
defparam \fifo_data~153 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][1] (
	.clk(clk),
	.d(\fifo_data~153_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~136 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~136_combout ),
	.cout());
defparam \fifo_data~136 .lut_mask = 16'hEEEE;
defparam \fifo_data~136 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][1] (
	.clk(clk),
	.d(\fifo_data~136_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~119 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~119_combout ),
	.cout());
defparam \fifo_data~119 .lut_mask = 16'hEEEE;
defparam \fifo_data~119 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][1] (
	.clk(clk),
	.d(\fifo_data~119_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~102 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~102_combout ),
	.cout());
defparam \fifo_data~102 .lut_mask = 16'hEEEE;
defparam \fifo_data~102 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][1] (
	.clk(clk),
	.d(\fifo_data~102_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~85 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~85_combout ),
	.cout());
defparam \fifo_data~85 .lut_mask = 16'hEEEE;
defparam \fifo_data~85 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][1] (
	.clk(clk),
	.d(\fifo_data~85_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~68 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~68_combout ),
	.cout());
defparam \fifo_data~68 .lut_mask = 16'hEEEE;
defparam \fifo_data~68 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][1] (
	.clk(clk),
	.d(\fifo_data~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~51 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~51_combout ),
	.cout());
defparam \fifo_data~51 .lut_mask = 16'hEEEE;
defparam \fifo_data~51 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][1] (
	.clk(clk),
	.d(\fifo_data~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~34 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~34_combout ),
	.cout());
defparam \fifo_data~34 .lut_mask = 16'hEEEE;
defparam \fifo_data~34 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][1] (
	.clk(clk),
	.d(\fifo_data~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~17 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~17_combout ),
	.cout());
defparam \fifo_data~17 .lut_mask = 16'hEEEE;
defparam \fifo_data~17 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][1] (
	.clk(clk),
	.d(\fifo_data~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][1] .power_up = "low";

cycloneive_lcell_comb \fifo_data~0 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~0_combout ),
	.cout());
defparam \fifo_data~0 .lut_mask = 16'hEEEE;
defparam \fifo_data~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~256 (
	.dataa(reset_n),
	.datab(Mux16),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~256_combout ),
	.cout());
defparam \fifo_data~256 .lut_mask = 16'hEEEE;
defparam \fifo_data~256 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\fifo_data~256_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~239 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~239_combout ),
	.cout());
defparam \fifo_data~239 .lut_mask = 16'hEEEE;
defparam \fifo_data~239 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][0] (
	.clk(clk),
	.d(\fifo_data~239_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~222 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~222_combout ),
	.cout());
defparam \fifo_data~222 .lut_mask = 16'hEEEE;
defparam \fifo_data~222 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][0] (
	.clk(clk),
	.d(\fifo_data~222_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~205 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~205_combout ),
	.cout());
defparam \fifo_data~205 .lut_mask = 16'hEEEE;
defparam \fifo_data~205 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][0] (
	.clk(clk),
	.d(\fifo_data~205_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~188 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~188_combout ),
	.cout());
defparam \fifo_data~188 .lut_mask = 16'hEEEE;
defparam \fifo_data~188 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][0] (
	.clk(clk),
	.d(\fifo_data~188_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~171 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~171_combout ),
	.cout());
defparam \fifo_data~171 .lut_mask = 16'hEEEE;
defparam \fifo_data~171 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][0] (
	.clk(clk),
	.d(\fifo_data~171_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~154 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~154_combout ),
	.cout());
defparam \fifo_data~154 .lut_mask = 16'hEEEE;
defparam \fifo_data~154 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][0] (
	.clk(clk),
	.d(\fifo_data~154_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~137 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~137_combout ),
	.cout());
defparam \fifo_data~137 .lut_mask = 16'hEEEE;
defparam \fifo_data~137 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][0] (
	.clk(clk),
	.d(\fifo_data~137_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~120 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~120_combout ),
	.cout());
defparam \fifo_data~120 .lut_mask = 16'hEEEE;
defparam \fifo_data~120 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][0] (
	.clk(clk),
	.d(\fifo_data~120_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~103 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~103_combout ),
	.cout());
defparam \fifo_data~103 .lut_mask = 16'hEEEE;
defparam \fifo_data~103 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][0] (
	.clk(clk),
	.d(\fifo_data~103_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~86 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~86_combout ),
	.cout());
defparam \fifo_data~86 .lut_mask = 16'hEEEE;
defparam \fifo_data~86 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][0] (
	.clk(clk),
	.d(\fifo_data~86_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~69 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~69_combout ),
	.cout());
defparam \fifo_data~69 .lut_mask = 16'hEEEE;
defparam \fifo_data~69 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][0] (
	.clk(clk),
	.d(\fifo_data~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~52 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~52_combout ),
	.cout());
defparam \fifo_data~52 .lut_mask = 16'hEEEE;
defparam \fifo_data~52 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][0] (
	.clk(clk),
	.d(\fifo_data~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~35 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~35_combout ),
	.cout());
defparam \fifo_data~35 .lut_mask = 16'hEEEE;
defparam \fifo_data~35 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][0] (
	.clk(clk),
	.d(\fifo_data~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~18 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~18_combout ),
	.cout());
defparam \fifo_data~18 .lut_mask = 16'hEEEE;
defparam \fifo_data~18 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][0] (
	.clk(clk),
	.d(\fifo_data~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][0] .power_up = "low";

cycloneive_lcell_comb \fifo_data~1 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~1_combout ),
	.cout());
defparam \fifo_data~1 .lut_mask = 16'hEEEE;
defparam \fifo_data~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~257 (
	.dataa(reset_n),
	.datab(Mux14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~257_combout ),
	.cout());
defparam \fifo_data~257 .lut_mask = 16'hEEEE;
defparam \fifo_data~257 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\fifo_data~257_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~240 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~240_combout ),
	.cout());
defparam \fifo_data~240 .lut_mask = 16'hEEEE;
defparam \fifo_data~240 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][2] (
	.clk(clk),
	.d(\fifo_data~240_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~223 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~223_combout ),
	.cout());
defparam \fifo_data~223 .lut_mask = 16'hEEEE;
defparam \fifo_data~223 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][2] (
	.clk(clk),
	.d(\fifo_data~223_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~206 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~206_combout ),
	.cout());
defparam \fifo_data~206 .lut_mask = 16'hEEEE;
defparam \fifo_data~206 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][2] (
	.clk(clk),
	.d(\fifo_data~206_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~189 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~189_combout ),
	.cout());
defparam \fifo_data~189 .lut_mask = 16'hEEEE;
defparam \fifo_data~189 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][2] (
	.clk(clk),
	.d(\fifo_data~189_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~172 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~172_combout ),
	.cout());
defparam \fifo_data~172 .lut_mask = 16'hEEEE;
defparam \fifo_data~172 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][2] (
	.clk(clk),
	.d(\fifo_data~172_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~155 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~155_combout ),
	.cout());
defparam \fifo_data~155 .lut_mask = 16'hEEEE;
defparam \fifo_data~155 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][2] (
	.clk(clk),
	.d(\fifo_data~155_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~138 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~138_combout ),
	.cout());
defparam \fifo_data~138 .lut_mask = 16'hEEEE;
defparam \fifo_data~138 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][2] (
	.clk(clk),
	.d(\fifo_data~138_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~121 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~121_combout ),
	.cout());
defparam \fifo_data~121 .lut_mask = 16'hEEEE;
defparam \fifo_data~121 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][2] (
	.clk(clk),
	.d(\fifo_data~121_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~104 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~104_combout ),
	.cout());
defparam \fifo_data~104 .lut_mask = 16'hEEEE;
defparam \fifo_data~104 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][2] (
	.clk(clk),
	.d(\fifo_data~104_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~87 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~87_combout ),
	.cout());
defparam \fifo_data~87 .lut_mask = 16'hEEEE;
defparam \fifo_data~87 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][2] (
	.clk(clk),
	.d(\fifo_data~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~70 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~70_combout ),
	.cout());
defparam \fifo_data~70 .lut_mask = 16'hEEEE;
defparam \fifo_data~70 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][2] (
	.clk(clk),
	.d(\fifo_data~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~53 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~53_combout ),
	.cout());
defparam \fifo_data~53 .lut_mask = 16'hEEEE;
defparam \fifo_data~53 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][2] (
	.clk(clk),
	.d(\fifo_data~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~36 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~36_combout ),
	.cout());
defparam \fifo_data~36 .lut_mask = 16'hEEEE;
defparam \fifo_data~36 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][2] (
	.clk(clk),
	.d(\fifo_data~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~19 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~19_combout ),
	.cout());
defparam \fifo_data~19 .lut_mask = 16'hEEEE;
defparam \fifo_data~19 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][2] (
	.clk(clk),
	.d(\fifo_data~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][2] .power_up = "low";

cycloneive_lcell_comb \fifo_data~2 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~2_combout ),
	.cout());
defparam \fifo_data~2 .lut_mask = 16'hEEEE;
defparam \fifo_data~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~258 (
	.dataa(reset_n),
	.datab(Mux13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~258_combout ),
	.cout());
defparam \fifo_data~258 .lut_mask = 16'hEEEE;
defparam \fifo_data~258 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\fifo_data~258_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~241 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~241_combout ),
	.cout());
defparam \fifo_data~241 .lut_mask = 16'hEEEE;
defparam \fifo_data~241 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][3] (
	.clk(clk),
	.d(\fifo_data~241_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~224 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~224_combout ),
	.cout());
defparam \fifo_data~224 .lut_mask = 16'hEEEE;
defparam \fifo_data~224 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][3] (
	.clk(clk),
	.d(\fifo_data~224_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~207 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~207_combout ),
	.cout());
defparam \fifo_data~207 .lut_mask = 16'hEEEE;
defparam \fifo_data~207 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][3] (
	.clk(clk),
	.d(\fifo_data~207_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~190 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~190_combout ),
	.cout());
defparam \fifo_data~190 .lut_mask = 16'hEEEE;
defparam \fifo_data~190 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][3] (
	.clk(clk),
	.d(\fifo_data~190_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~173 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~173_combout ),
	.cout());
defparam \fifo_data~173 .lut_mask = 16'hEEEE;
defparam \fifo_data~173 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][3] (
	.clk(clk),
	.d(\fifo_data~173_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~156 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~156_combout ),
	.cout());
defparam \fifo_data~156 .lut_mask = 16'hEEEE;
defparam \fifo_data~156 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][3] (
	.clk(clk),
	.d(\fifo_data~156_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~139 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~139_combout ),
	.cout());
defparam \fifo_data~139 .lut_mask = 16'hEEEE;
defparam \fifo_data~139 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][3] (
	.clk(clk),
	.d(\fifo_data~139_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~122 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~122_combout ),
	.cout());
defparam \fifo_data~122 .lut_mask = 16'hEEEE;
defparam \fifo_data~122 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][3] (
	.clk(clk),
	.d(\fifo_data~122_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~105 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~105_combout ),
	.cout());
defparam \fifo_data~105 .lut_mask = 16'hEEEE;
defparam \fifo_data~105 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][3] (
	.clk(clk),
	.d(\fifo_data~105_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~88 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~88_combout ),
	.cout());
defparam \fifo_data~88 .lut_mask = 16'hEEEE;
defparam \fifo_data~88 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][3] (
	.clk(clk),
	.d(\fifo_data~88_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~71 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~71_combout ),
	.cout());
defparam \fifo_data~71 .lut_mask = 16'hEEEE;
defparam \fifo_data~71 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][3] (
	.clk(clk),
	.d(\fifo_data~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~54 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~54_combout ),
	.cout());
defparam \fifo_data~54 .lut_mask = 16'hEEEE;
defparam \fifo_data~54 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][3] (
	.clk(clk),
	.d(\fifo_data~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~37 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~37_combout ),
	.cout());
defparam \fifo_data~37 .lut_mask = 16'hEEEE;
defparam \fifo_data~37 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][3] (
	.clk(clk),
	.d(\fifo_data~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~20 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~20_combout ),
	.cout());
defparam \fifo_data~20 .lut_mask = 16'hEEEE;
defparam \fifo_data~20 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][3] (
	.clk(clk),
	.d(\fifo_data~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][3] .power_up = "low";

cycloneive_lcell_comb \fifo_data~3 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~3_combout ),
	.cout());
defparam \fifo_data~3 .lut_mask = 16'hEEEE;
defparam \fifo_data~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~259 (
	.dataa(reset_n),
	.datab(Mux12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~259_combout ),
	.cout());
defparam \fifo_data~259 .lut_mask = 16'hEEEE;
defparam \fifo_data~259 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\fifo_data~259_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~242 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~242_combout ),
	.cout());
defparam \fifo_data~242 .lut_mask = 16'hEEEE;
defparam \fifo_data~242 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][4] (
	.clk(clk),
	.d(\fifo_data~242_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~225 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~225_combout ),
	.cout());
defparam \fifo_data~225 .lut_mask = 16'hEEEE;
defparam \fifo_data~225 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][4] (
	.clk(clk),
	.d(\fifo_data~225_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~208 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~208_combout ),
	.cout());
defparam \fifo_data~208 .lut_mask = 16'hEEEE;
defparam \fifo_data~208 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][4] (
	.clk(clk),
	.d(\fifo_data~208_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~191 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~191_combout ),
	.cout());
defparam \fifo_data~191 .lut_mask = 16'hEEEE;
defparam \fifo_data~191 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][4] (
	.clk(clk),
	.d(\fifo_data~191_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~174 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~174_combout ),
	.cout());
defparam \fifo_data~174 .lut_mask = 16'hEEEE;
defparam \fifo_data~174 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][4] (
	.clk(clk),
	.d(\fifo_data~174_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~157 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~157_combout ),
	.cout());
defparam \fifo_data~157 .lut_mask = 16'hEEEE;
defparam \fifo_data~157 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][4] (
	.clk(clk),
	.d(\fifo_data~157_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~140 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~140_combout ),
	.cout());
defparam \fifo_data~140 .lut_mask = 16'hEEEE;
defparam \fifo_data~140 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][4] (
	.clk(clk),
	.d(\fifo_data~140_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~123 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~123_combout ),
	.cout());
defparam \fifo_data~123 .lut_mask = 16'hEEEE;
defparam \fifo_data~123 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][4] (
	.clk(clk),
	.d(\fifo_data~123_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~106 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~106_combout ),
	.cout());
defparam \fifo_data~106 .lut_mask = 16'hEEEE;
defparam \fifo_data~106 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][4] (
	.clk(clk),
	.d(\fifo_data~106_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~89 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~89_combout ),
	.cout());
defparam \fifo_data~89 .lut_mask = 16'hEEEE;
defparam \fifo_data~89 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][4] (
	.clk(clk),
	.d(\fifo_data~89_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~72 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~72_combout ),
	.cout());
defparam \fifo_data~72 .lut_mask = 16'hEEEE;
defparam \fifo_data~72 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][4] (
	.clk(clk),
	.d(\fifo_data~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~55 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~55_combout ),
	.cout());
defparam \fifo_data~55 .lut_mask = 16'hEEEE;
defparam \fifo_data~55 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][4] (
	.clk(clk),
	.d(\fifo_data~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~38 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~38_combout ),
	.cout());
defparam \fifo_data~38 .lut_mask = 16'hEEEE;
defparam \fifo_data~38 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][4] (
	.clk(clk),
	.d(\fifo_data~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~21 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~21_combout ),
	.cout());
defparam \fifo_data~21 .lut_mask = 16'hEEEE;
defparam \fifo_data~21 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][4] (
	.clk(clk),
	.d(\fifo_data~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][4] .power_up = "low";

cycloneive_lcell_comb \fifo_data~4 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~4_combout ),
	.cout());
defparam \fifo_data~4 .lut_mask = 16'hEEEE;
defparam \fifo_data~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~260 (
	.dataa(reset_n),
	.datab(Mux11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~260_combout ),
	.cout());
defparam \fifo_data~260 .lut_mask = 16'hEEEE;
defparam \fifo_data~260 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\fifo_data~260_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~243 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~243_combout ),
	.cout());
defparam \fifo_data~243 .lut_mask = 16'hEEEE;
defparam \fifo_data~243 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][5] (
	.clk(clk),
	.d(\fifo_data~243_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~226 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~226_combout ),
	.cout());
defparam \fifo_data~226 .lut_mask = 16'hEEEE;
defparam \fifo_data~226 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][5] (
	.clk(clk),
	.d(\fifo_data~226_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~209 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~209_combout ),
	.cout());
defparam \fifo_data~209 .lut_mask = 16'hEEEE;
defparam \fifo_data~209 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][5] (
	.clk(clk),
	.d(\fifo_data~209_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~192 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~192_combout ),
	.cout());
defparam \fifo_data~192 .lut_mask = 16'hEEEE;
defparam \fifo_data~192 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][5] (
	.clk(clk),
	.d(\fifo_data~192_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~175 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~175_combout ),
	.cout());
defparam \fifo_data~175 .lut_mask = 16'hEEEE;
defparam \fifo_data~175 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][5] (
	.clk(clk),
	.d(\fifo_data~175_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~158 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~158_combout ),
	.cout());
defparam \fifo_data~158 .lut_mask = 16'hEEEE;
defparam \fifo_data~158 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][5] (
	.clk(clk),
	.d(\fifo_data~158_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~141 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~141_combout ),
	.cout());
defparam \fifo_data~141 .lut_mask = 16'hEEEE;
defparam \fifo_data~141 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][5] (
	.clk(clk),
	.d(\fifo_data~141_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~124 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~124_combout ),
	.cout());
defparam \fifo_data~124 .lut_mask = 16'hEEEE;
defparam \fifo_data~124 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][5] (
	.clk(clk),
	.d(\fifo_data~124_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~107 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~107_combout ),
	.cout());
defparam \fifo_data~107 .lut_mask = 16'hEEEE;
defparam \fifo_data~107 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][5] (
	.clk(clk),
	.d(\fifo_data~107_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~90 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~90_combout ),
	.cout());
defparam \fifo_data~90 .lut_mask = 16'hEEEE;
defparam \fifo_data~90 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][5] (
	.clk(clk),
	.d(\fifo_data~90_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~73 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~73_combout ),
	.cout());
defparam \fifo_data~73 .lut_mask = 16'hEEEE;
defparam \fifo_data~73 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][5] (
	.clk(clk),
	.d(\fifo_data~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~56 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~56_combout ),
	.cout());
defparam \fifo_data~56 .lut_mask = 16'hEEEE;
defparam \fifo_data~56 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][5] (
	.clk(clk),
	.d(\fifo_data~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~39 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~39_combout ),
	.cout());
defparam \fifo_data~39 .lut_mask = 16'hEEEE;
defparam \fifo_data~39 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][5] (
	.clk(clk),
	.d(\fifo_data~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~22 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~22_combout ),
	.cout());
defparam \fifo_data~22 .lut_mask = 16'hEEEE;
defparam \fifo_data~22 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][5] (
	.clk(clk),
	.d(\fifo_data~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][5]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][5] .power_up = "low";

cycloneive_lcell_comb \fifo_data~5 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~5_combout ),
	.cout());
defparam \fifo_data~5 .lut_mask = 16'hEEEE;
defparam \fifo_data~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~261 (
	.dataa(reset_n),
	.datab(Mux10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~261_combout ),
	.cout());
defparam \fifo_data~261 .lut_mask = 16'hEEEE;
defparam \fifo_data~261 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\fifo_data~261_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~244 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~244_combout ),
	.cout());
defparam \fifo_data~244 .lut_mask = 16'hEEEE;
defparam \fifo_data~244 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][6] (
	.clk(clk),
	.d(\fifo_data~244_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~227 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~227_combout ),
	.cout());
defparam \fifo_data~227 .lut_mask = 16'hEEEE;
defparam \fifo_data~227 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][6] (
	.clk(clk),
	.d(\fifo_data~227_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~210 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~210_combout ),
	.cout());
defparam \fifo_data~210 .lut_mask = 16'hEEEE;
defparam \fifo_data~210 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][6] (
	.clk(clk),
	.d(\fifo_data~210_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~193 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~193_combout ),
	.cout());
defparam \fifo_data~193 .lut_mask = 16'hEEEE;
defparam \fifo_data~193 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][6] (
	.clk(clk),
	.d(\fifo_data~193_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~176 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~176_combout ),
	.cout());
defparam \fifo_data~176 .lut_mask = 16'hEEEE;
defparam \fifo_data~176 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][6] (
	.clk(clk),
	.d(\fifo_data~176_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~159 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~159_combout ),
	.cout());
defparam \fifo_data~159 .lut_mask = 16'hEEEE;
defparam \fifo_data~159 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][6] (
	.clk(clk),
	.d(\fifo_data~159_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~142 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~142_combout ),
	.cout());
defparam \fifo_data~142 .lut_mask = 16'hEEEE;
defparam \fifo_data~142 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][6] (
	.clk(clk),
	.d(\fifo_data~142_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~125 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~125_combout ),
	.cout());
defparam \fifo_data~125 .lut_mask = 16'hEEEE;
defparam \fifo_data~125 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][6] (
	.clk(clk),
	.d(\fifo_data~125_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~108 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~108_combout ),
	.cout());
defparam \fifo_data~108 .lut_mask = 16'hEEEE;
defparam \fifo_data~108 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][6] (
	.clk(clk),
	.d(\fifo_data~108_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~91 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~91_combout ),
	.cout());
defparam \fifo_data~91 .lut_mask = 16'hEEEE;
defparam \fifo_data~91 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][6] (
	.clk(clk),
	.d(\fifo_data~91_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~74 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~74_combout ),
	.cout());
defparam \fifo_data~74 .lut_mask = 16'hEEEE;
defparam \fifo_data~74 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][6] (
	.clk(clk),
	.d(\fifo_data~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~57 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~57_combout ),
	.cout());
defparam \fifo_data~57 .lut_mask = 16'hEEEE;
defparam \fifo_data~57 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][6] (
	.clk(clk),
	.d(\fifo_data~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~40 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~40_combout ),
	.cout());
defparam \fifo_data~40 .lut_mask = 16'hEEEE;
defparam \fifo_data~40 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][6] (
	.clk(clk),
	.d(\fifo_data~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~23 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~23_combout ),
	.cout());
defparam \fifo_data~23 .lut_mask = 16'hEEEE;
defparam \fifo_data~23 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][6] (
	.clk(clk),
	.d(\fifo_data~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][6]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][6] .power_up = "low";

cycloneive_lcell_comb \fifo_data~6 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~6_combout ),
	.cout());
defparam \fifo_data~6 .lut_mask = 16'hEEEE;
defparam \fifo_data~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~262 (
	.dataa(reset_n),
	.datab(Mux9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~262_combout ),
	.cout());
defparam \fifo_data~262 .lut_mask = 16'hEEEE;
defparam \fifo_data~262 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\fifo_data~262_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~245 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~245_combout ),
	.cout());
defparam \fifo_data~245 .lut_mask = 16'hEEEE;
defparam \fifo_data~245 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][7] (
	.clk(clk),
	.d(\fifo_data~245_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~228 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~228_combout ),
	.cout());
defparam \fifo_data~228 .lut_mask = 16'hEEEE;
defparam \fifo_data~228 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][7] (
	.clk(clk),
	.d(\fifo_data~228_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~211 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~211_combout ),
	.cout());
defparam \fifo_data~211 .lut_mask = 16'hEEEE;
defparam \fifo_data~211 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][7] (
	.clk(clk),
	.d(\fifo_data~211_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~194 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~194_combout ),
	.cout());
defparam \fifo_data~194 .lut_mask = 16'hEEEE;
defparam \fifo_data~194 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][7] (
	.clk(clk),
	.d(\fifo_data~194_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~177 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~177_combout ),
	.cout());
defparam \fifo_data~177 .lut_mask = 16'hEEEE;
defparam \fifo_data~177 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][7] (
	.clk(clk),
	.d(\fifo_data~177_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~160 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~160_combout ),
	.cout());
defparam \fifo_data~160 .lut_mask = 16'hEEEE;
defparam \fifo_data~160 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][7] (
	.clk(clk),
	.d(\fifo_data~160_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~143 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~143_combout ),
	.cout());
defparam \fifo_data~143 .lut_mask = 16'hEEEE;
defparam \fifo_data~143 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][7] (
	.clk(clk),
	.d(\fifo_data~143_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~126 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~126_combout ),
	.cout());
defparam \fifo_data~126 .lut_mask = 16'hEEEE;
defparam \fifo_data~126 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][7] (
	.clk(clk),
	.d(\fifo_data~126_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~109 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~109_combout ),
	.cout());
defparam \fifo_data~109 .lut_mask = 16'hEEEE;
defparam \fifo_data~109 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][7] (
	.clk(clk),
	.d(\fifo_data~109_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~92 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~92_combout ),
	.cout());
defparam \fifo_data~92 .lut_mask = 16'hEEEE;
defparam \fifo_data~92 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][7] (
	.clk(clk),
	.d(\fifo_data~92_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~75 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~75_combout ),
	.cout());
defparam \fifo_data~75 .lut_mask = 16'hEEEE;
defparam \fifo_data~75 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][7] (
	.clk(clk),
	.d(\fifo_data~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~58 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~58_combout ),
	.cout());
defparam \fifo_data~58 .lut_mask = 16'hEEEE;
defparam \fifo_data~58 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][7] (
	.clk(clk),
	.d(\fifo_data~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~41 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~41_combout ),
	.cout());
defparam \fifo_data~41 .lut_mask = 16'hEEEE;
defparam \fifo_data~41 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][7] (
	.clk(clk),
	.d(\fifo_data~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~24 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~24_combout ),
	.cout());
defparam \fifo_data~24 .lut_mask = 16'hEEEE;
defparam \fifo_data~24 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][7] (
	.clk(clk),
	.d(\fifo_data~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][7]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][7] .power_up = "low";

cycloneive_lcell_comb \fifo_data~7 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~7_combout ),
	.cout());
defparam \fifo_data~7 .lut_mask = 16'hEEEE;
defparam \fifo_data~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~263 (
	.dataa(reset_n),
	.datab(Mux8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~263_combout ),
	.cout());
defparam \fifo_data~263 .lut_mask = 16'hEEEE;
defparam \fifo_data~263 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\fifo_data~263_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~246 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~246_combout ),
	.cout());
defparam \fifo_data~246 .lut_mask = 16'hEEEE;
defparam \fifo_data~246 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][8] (
	.clk(clk),
	.d(\fifo_data~246_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~229 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~229_combout ),
	.cout());
defparam \fifo_data~229 .lut_mask = 16'hEEEE;
defparam \fifo_data~229 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][8] (
	.clk(clk),
	.d(\fifo_data~229_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~212 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~212_combout ),
	.cout());
defparam \fifo_data~212 .lut_mask = 16'hEEEE;
defparam \fifo_data~212 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][8] (
	.clk(clk),
	.d(\fifo_data~212_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~195 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~195_combout ),
	.cout());
defparam \fifo_data~195 .lut_mask = 16'hEEEE;
defparam \fifo_data~195 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][8] (
	.clk(clk),
	.d(\fifo_data~195_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~178 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~178_combout ),
	.cout());
defparam \fifo_data~178 .lut_mask = 16'hEEEE;
defparam \fifo_data~178 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][8] (
	.clk(clk),
	.d(\fifo_data~178_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~161 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~161_combout ),
	.cout());
defparam \fifo_data~161 .lut_mask = 16'hEEEE;
defparam \fifo_data~161 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][8] (
	.clk(clk),
	.d(\fifo_data~161_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~144 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~144_combout ),
	.cout());
defparam \fifo_data~144 .lut_mask = 16'hEEEE;
defparam \fifo_data~144 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][8] (
	.clk(clk),
	.d(\fifo_data~144_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~127 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~127_combout ),
	.cout());
defparam \fifo_data~127 .lut_mask = 16'hEEEE;
defparam \fifo_data~127 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][8] (
	.clk(clk),
	.d(\fifo_data~127_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~110 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~110_combout ),
	.cout());
defparam \fifo_data~110 .lut_mask = 16'hEEEE;
defparam \fifo_data~110 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][8] (
	.clk(clk),
	.d(\fifo_data~110_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~93 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~93_combout ),
	.cout());
defparam \fifo_data~93 .lut_mask = 16'hEEEE;
defparam \fifo_data~93 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][8] (
	.clk(clk),
	.d(\fifo_data~93_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~76 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~76_combout ),
	.cout());
defparam \fifo_data~76 .lut_mask = 16'hEEEE;
defparam \fifo_data~76 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][8] (
	.clk(clk),
	.d(\fifo_data~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~59 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~59_combout ),
	.cout());
defparam \fifo_data~59 .lut_mask = 16'hEEEE;
defparam \fifo_data~59 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][8] (
	.clk(clk),
	.d(\fifo_data~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~42 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~42_combout ),
	.cout());
defparam \fifo_data~42 .lut_mask = 16'hEEEE;
defparam \fifo_data~42 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][8] (
	.clk(clk),
	.d(\fifo_data~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~25 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~25_combout ),
	.cout());
defparam \fifo_data~25 .lut_mask = 16'hEEEE;
defparam \fifo_data~25 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][8] (
	.clk(clk),
	.d(\fifo_data~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][8]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][8] .power_up = "low";

cycloneive_lcell_comb \fifo_data~8 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~8_combout ),
	.cout());
defparam \fifo_data~8 .lut_mask = 16'hEEEE;
defparam \fifo_data~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~264 (
	.dataa(reset_n),
	.datab(Mux7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~264_combout ),
	.cout());
defparam \fifo_data~264 .lut_mask = 16'hEEEE;
defparam \fifo_data~264 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\fifo_data~264_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~247 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~247_combout ),
	.cout());
defparam \fifo_data~247 .lut_mask = 16'hEEEE;
defparam \fifo_data~247 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][9] (
	.clk(clk),
	.d(\fifo_data~247_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~230 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~230_combout ),
	.cout());
defparam \fifo_data~230 .lut_mask = 16'hEEEE;
defparam \fifo_data~230 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][9] (
	.clk(clk),
	.d(\fifo_data~230_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~213 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~213_combout ),
	.cout());
defparam \fifo_data~213 .lut_mask = 16'hEEEE;
defparam \fifo_data~213 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][9] (
	.clk(clk),
	.d(\fifo_data~213_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~196 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~196_combout ),
	.cout());
defparam \fifo_data~196 .lut_mask = 16'hEEEE;
defparam \fifo_data~196 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][9] (
	.clk(clk),
	.d(\fifo_data~196_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~179 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~179_combout ),
	.cout());
defparam \fifo_data~179 .lut_mask = 16'hEEEE;
defparam \fifo_data~179 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][9] (
	.clk(clk),
	.d(\fifo_data~179_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~162 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~162_combout ),
	.cout());
defparam \fifo_data~162 .lut_mask = 16'hEEEE;
defparam \fifo_data~162 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][9] (
	.clk(clk),
	.d(\fifo_data~162_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~145 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~145_combout ),
	.cout());
defparam \fifo_data~145 .lut_mask = 16'hEEEE;
defparam \fifo_data~145 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][9] (
	.clk(clk),
	.d(\fifo_data~145_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~128 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~128_combout ),
	.cout());
defparam \fifo_data~128 .lut_mask = 16'hEEEE;
defparam \fifo_data~128 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][9] (
	.clk(clk),
	.d(\fifo_data~128_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~111 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~111_combout ),
	.cout());
defparam \fifo_data~111 .lut_mask = 16'hEEEE;
defparam \fifo_data~111 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][9] (
	.clk(clk),
	.d(\fifo_data~111_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~94 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~94_combout ),
	.cout());
defparam \fifo_data~94 .lut_mask = 16'hEEEE;
defparam \fifo_data~94 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][9] (
	.clk(clk),
	.d(\fifo_data~94_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~77 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~77_combout ),
	.cout());
defparam \fifo_data~77 .lut_mask = 16'hEEEE;
defparam \fifo_data~77 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][9] (
	.clk(clk),
	.d(\fifo_data~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~60 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~60_combout ),
	.cout());
defparam \fifo_data~60 .lut_mask = 16'hEEEE;
defparam \fifo_data~60 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][9] (
	.clk(clk),
	.d(\fifo_data~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~43 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~43_combout ),
	.cout());
defparam \fifo_data~43 .lut_mask = 16'hEEEE;
defparam \fifo_data~43 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][9] (
	.clk(clk),
	.d(\fifo_data~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~26 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~26_combout ),
	.cout());
defparam \fifo_data~26 .lut_mask = 16'hEEEE;
defparam \fifo_data~26 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][9] (
	.clk(clk),
	.d(\fifo_data~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][9]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][9] .power_up = "low";

cycloneive_lcell_comb \fifo_data~9 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~9_combout ),
	.cout());
defparam \fifo_data~9 .lut_mask = 16'hEEEE;
defparam \fifo_data~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~265 (
	.dataa(reset_n),
	.datab(Mux6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~265_combout ),
	.cout());
defparam \fifo_data~265 .lut_mask = 16'hEEEE;
defparam \fifo_data~265 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\fifo_data~265_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~248 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~248_combout ),
	.cout());
defparam \fifo_data~248 .lut_mask = 16'hEEEE;
defparam \fifo_data~248 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][10] (
	.clk(clk),
	.d(\fifo_data~248_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~231 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~231_combout ),
	.cout());
defparam \fifo_data~231 .lut_mask = 16'hEEEE;
defparam \fifo_data~231 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][10] (
	.clk(clk),
	.d(\fifo_data~231_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~214 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~214_combout ),
	.cout());
defparam \fifo_data~214 .lut_mask = 16'hEEEE;
defparam \fifo_data~214 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][10] (
	.clk(clk),
	.d(\fifo_data~214_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~197 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~197_combout ),
	.cout());
defparam \fifo_data~197 .lut_mask = 16'hEEEE;
defparam \fifo_data~197 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][10] (
	.clk(clk),
	.d(\fifo_data~197_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~180 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~180_combout ),
	.cout());
defparam \fifo_data~180 .lut_mask = 16'hEEEE;
defparam \fifo_data~180 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][10] (
	.clk(clk),
	.d(\fifo_data~180_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~163 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~163_combout ),
	.cout());
defparam \fifo_data~163 .lut_mask = 16'hEEEE;
defparam \fifo_data~163 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][10] (
	.clk(clk),
	.d(\fifo_data~163_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~146 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~146_combout ),
	.cout());
defparam \fifo_data~146 .lut_mask = 16'hEEEE;
defparam \fifo_data~146 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][10] (
	.clk(clk),
	.d(\fifo_data~146_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~129 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~129_combout ),
	.cout());
defparam \fifo_data~129 .lut_mask = 16'hEEEE;
defparam \fifo_data~129 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][10] (
	.clk(clk),
	.d(\fifo_data~129_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~112 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~112_combout ),
	.cout());
defparam \fifo_data~112 .lut_mask = 16'hEEEE;
defparam \fifo_data~112 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][10] (
	.clk(clk),
	.d(\fifo_data~112_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~95 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~95_combout ),
	.cout());
defparam \fifo_data~95 .lut_mask = 16'hEEEE;
defparam \fifo_data~95 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][10] (
	.clk(clk),
	.d(\fifo_data~95_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~78 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~78_combout ),
	.cout());
defparam \fifo_data~78 .lut_mask = 16'hEEEE;
defparam \fifo_data~78 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][10] (
	.clk(clk),
	.d(\fifo_data~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~61 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~61_combout ),
	.cout());
defparam \fifo_data~61 .lut_mask = 16'hEEEE;
defparam \fifo_data~61 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][10] (
	.clk(clk),
	.d(\fifo_data~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~44 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~44_combout ),
	.cout());
defparam \fifo_data~44 .lut_mask = 16'hEEEE;
defparam \fifo_data~44 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][10] (
	.clk(clk),
	.d(\fifo_data~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~27 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~27_combout ),
	.cout());
defparam \fifo_data~27 .lut_mask = 16'hEEEE;
defparam \fifo_data~27 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][10] (
	.clk(clk),
	.d(\fifo_data~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][10]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][10] .power_up = "low";

cycloneive_lcell_comb \fifo_data~10 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~10_combout ),
	.cout());
defparam \fifo_data~10 .lut_mask = 16'hEEEE;
defparam \fifo_data~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~266 (
	.dataa(reset_n),
	.datab(Mux5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~266_combout ),
	.cout());
defparam \fifo_data~266 .lut_mask = 16'hEEEE;
defparam \fifo_data~266 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\fifo_data~266_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~249 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~249_combout ),
	.cout());
defparam \fifo_data~249 .lut_mask = 16'hEEEE;
defparam \fifo_data~249 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][11] (
	.clk(clk),
	.d(\fifo_data~249_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~232 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~232_combout ),
	.cout());
defparam \fifo_data~232 .lut_mask = 16'hEEEE;
defparam \fifo_data~232 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][11] (
	.clk(clk),
	.d(\fifo_data~232_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~215 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~215_combout ),
	.cout());
defparam \fifo_data~215 .lut_mask = 16'hEEEE;
defparam \fifo_data~215 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][11] (
	.clk(clk),
	.d(\fifo_data~215_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~198 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~198_combout ),
	.cout());
defparam \fifo_data~198 .lut_mask = 16'hEEEE;
defparam \fifo_data~198 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][11] (
	.clk(clk),
	.d(\fifo_data~198_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~181 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~181_combout ),
	.cout());
defparam \fifo_data~181 .lut_mask = 16'hEEEE;
defparam \fifo_data~181 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][11] (
	.clk(clk),
	.d(\fifo_data~181_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~164 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~164_combout ),
	.cout());
defparam \fifo_data~164 .lut_mask = 16'hEEEE;
defparam \fifo_data~164 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][11] (
	.clk(clk),
	.d(\fifo_data~164_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~147 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~147_combout ),
	.cout());
defparam \fifo_data~147 .lut_mask = 16'hEEEE;
defparam \fifo_data~147 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][11] (
	.clk(clk),
	.d(\fifo_data~147_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~130 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~130_combout ),
	.cout());
defparam \fifo_data~130 .lut_mask = 16'hEEEE;
defparam \fifo_data~130 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][11] (
	.clk(clk),
	.d(\fifo_data~130_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~113 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~113_combout ),
	.cout());
defparam \fifo_data~113 .lut_mask = 16'hEEEE;
defparam \fifo_data~113 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][11] (
	.clk(clk),
	.d(\fifo_data~113_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~96 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~96_combout ),
	.cout());
defparam \fifo_data~96 .lut_mask = 16'hEEEE;
defparam \fifo_data~96 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][11] (
	.clk(clk),
	.d(\fifo_data~96_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~79 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~79_combout ),
	.cout());
defparam \fifo_data~79 .lut_mask = 16'hEEEE;
defparam \fifo_data~79 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][11] (
	.clk(clk),
	.d(\fifo_data~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~62 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~62_combout ),
	.cout());
defparam \fifo_data~62 .lut_mask = 16'hEEEE;
defparam \fifo_data~62 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][11] (
	.clk(clk),
	.d(\fifo_data~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~45 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~45_combout ),
	.cout());
defparam \fifo_data~45 .lut_mask = 16'hEEEE;
defparam \fifo_data~45 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][11] (
	.clk(clk),
	.d(\fifo_data~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~28 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~28_combout ),
	.cout());
defparam \fifo_data~28 .lut_mask = 16'hEEEE;
defparam \fifo_data~28 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][11] (
	.clk(clk),
	.d(\fifo_data~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][11]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][11] .power_up = "low";

cycloneive_lcell_comb \fifo_data~11 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~11_combout ),
	.cout());
defparam \fifo_data~11 .lut_mask = 16'hEEEE;
defparam \fifo_data~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~267 (
	.dataa(reset_n),
	.datab(Mux4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~267_combout ),
	.cout());
defparam \fifo_data~267 .lut_mask = 16'hEEEE;
defparam \fifo_data~267 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\fifo_data~267_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~250 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~250_combout ),
	.cout());
defparam \fifo_data~250 .lut_mask = 16'hEEEE;
defparam \fifo_data~250 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][12] (
	.clk(clk),
	.d(\fifo_data~250_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~233 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~233_combout ),
	.cout());
defparam \fifo_data~233 .lut_mask = 16'hEEEE;
defparam \fifo_data~233 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][12] (
	.clk(clk),
	.d(\fifo_data~233_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~216 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~216_combout ),
	.cout());
defparam \fifo_data~216 .lut_mask = 16'hEEEE;
defparam \fifo_data~216 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][12] (
	.clk(clk),
	.d(\fifo_data~216_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~199 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~199_combout ),
	.cout());
defparam \fifo_data~199 .lut_mask = 16'hEEEE;
defparam \fifo_data~199 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][12] (
	.clk(clk),
	.d(\fifo_data~199_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~182 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~182_combout ),
	.cout());
defparam \fifo_data~182 .lut_mask = 16'hEEEE;
defparam \fifo_data~182 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][12] (
	.clk(clk),
	.d(\fifo_data~182_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~165 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~165_combout ),
	.cout());
defparam \fifo_data~165 .lut_mask = 16'hEEEE;
defparam \fifo_data~165 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][12] (
	.clk(clk),
	.d(\fifo_data~165_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~148 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~148_combout ),
	.cout());
defparam \fifo_data~148 .lut_mask = 16'hEEEE;
defparam \fifo_data~148 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][12] (
	.clk(clk),
	.d(\fifo_data~148_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~131 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~131_combout ),
	.cout());
defparam \fifo_data~131 .lut_mask = 16'hEEEE;
defparam \fifo_data~131 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][12] (
	.clk(clk),
	.d(\fifo_data~131_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~114 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~114_combout ),
	.cout());
defparam \fifo_data~114 .lut_mask = 16'hEEEE;
defparam \fifo_data~114 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][12] (
	.clk(clk),
	.d(\fifo_data~114_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~97 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~97_combout ),
	.cout());
defparam \fifo_data~97 .lut_mask = 16'hEEEE;
defparam \fifo_data~97 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][12] (
	.clk(clk),
	.d(\fifo_data~97_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~80 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~80_combout ),
	.cout());
defparam \fifo_data~80 .lut_mask = 16'hEEEE;
defparam \fifo_data~80 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][12] (
	.clk(clk),
	.d(\fifo_data~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~63 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~63_combout ),
	.cout());
defparam \fifo_data~63 .lut_mask = 16'hEEEE;
defparam \fifo_data~63 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][12] (
	.clk(clk),
	.d(\fifo_data~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~46 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~46_combout ),
	.cout());
defparam \fifo_data~46 .lut_mask = 16'hEEEE;
defparam \fifo_data~46 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][12] (
	.clk(clk),
	.d(\fifo_data~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~29 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~29_combout ),
	.cout());
defparam \fifo_data~29 .lut_mask = 16'hEEEE;
defparam \fifo_data~29 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][12] (
	.clk(clk),
	.d(\fifo_data~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][12]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][12] .power_up = "low";

cycloneive_lcell_comb \fifo_data~12 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~12_combout ),
	.cout());
defparam \fifo_data~12 .lut_mask = 16'hEEEE;
defparam \fifo_data~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~268 (
	.dataa(reset_n),
	.datab(Mux3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~268_combout ),
	.cout());
defparam \fifo_data~268 .lut_mask = 16'hEEEE;
defparam \fifo_data~268 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\fifo_data~268_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~251 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~251_combout ),
	.cout());
defparam \fifo_data~251 .lut_mask = 16'hEEEE;
defparam \fifo_data~251 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][13] (
	.clk(clk),
	.d(\fifo_data~251_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~234 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~234_combout ),
	.cout());
defparam \fifo_data~234 .lut_mask = 16'hEEEE;
defparam \fifo_data~234 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][13] (
	.clk(clk),
	.d(\fifo_data~234_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~217 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~217_combout ),
	.cout());
defparam \fifo_data~217 .lut_mask = 16'hEEEE;
defparam \fifo_data~217 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][13] (
	.clk(clk),
	.d(\fifo_data~217_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~200 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~200_combout ),
	.cout());
defparam \fifo_data~200 .lut_mask = 16'hEEEE;
defparam \fifo_data~200 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][13] (
	.clk(clk),
	.d(\fifo_data~200_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~183 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~183_combout ),
	.cout());
defparam \fifo_data~183 .lut_mask = 16'hEEEE;
defparam \fifo_data~183 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][13] (
	.clk(clk),
	.d(\fifo_data~183_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~166 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~166_combout ),
	.cout());
defparam \fifo_data~166 .lut_mask = 16'hEEEE;
defparam \fifo_data~166 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][13] (
	.clk(clk),
	.d(\fifo_data~166_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~149 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~149_combout ),
	.cout());
defparam \fifo_data~149 .lut_mask = 16'hEEEE;
defparam \fifo_data~149 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][13] (
	.clk(clk),
	.d(\fifo_data~149_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~132 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~132_combout ),
	.cout());
defparam \fifo_data~132 .lut_mask = 16'hEEEE;
defparam \fifo_data~132 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][13] (
	.clk(clk),
	.d(\fifo_data~132_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~115 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~115_combout ),
	.cout());
defparam \fifo_data~115 .lut_mask = 16'hEEEE;
defparam \fifo_data~115 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][13] (
	.clk(clk),
	.d(\fifo_data~115_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~98 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~98_combout ),
	.cout());
defparam \fifo_data~98 .lut_mask = 16'hEEEE;
defparam \fifo_data~98 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][13] (
	.clk(clk),
	.d(\fifo_data~98_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~81 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~81_combout ),
	.cout());
defparam \fifo_data~81 .lut_mask = 16'hEEEE;
defparam \fifo_data~81 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][13] (
	.clk(clk),
	.d(\fifo_data~81_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~64 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~64_combout ),
	.cout());
defparam \fifo_data~64 .lut_mask = 16'hEEEE;
defparam \fifo_data~64 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][13] (
	.clk(clk),
	.d(\fifo_data~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~47 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~47_combout ),
	.cout());
defparam \fifo_data~47 .lut_mask = 16'hEEEE;
defparam \fifo_data~47 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][13] (
	.clk(clk),
	.d(\fifo_data~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~30 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~30_combout ),
	.cout());
defparam \fifo_data~30 .lut_mask = 16'hEEEE;
defparam \fifo_data~30 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][13] (
	.clk(clk),
	.d(\fifo_data~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][13]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][13] .power_up = "low";

cycloneive_lcell_comb \fifo_data~13 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~13_combout ),
	.cout());
defparam \fifo_data~13 .lut_mask = 16'hEEEE;
defparam \fifo_data~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~269 (
	.dataa(reset_n),
	.datab(Mux2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~269_combout ),
	.cout());
defparam \fifo_data~269 .lut_mask = 16'hEEEE;
defparam \fifo_data~269 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\fifo_data~269_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~252 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~252_combout ),
	.cout());
defparam \fifo_data~252 .lut_mask = 16'hEEEE;
defparam \fifo_data~252 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][14] (
	.clk(clk),
	.d(\fifo_data~252_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~235 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~235_combout ),
	.cout());
defparam \fifo_data~235 .lut_mask = 16'hEEEE;
defparam \fifo_data~235 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][14] (
	.clk(clk),
	.d(\fifo_data~235_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~218 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~218_combout ),
	.cout());
defparam \fifo_data~218 .lut_mask = 16'hEEEE;
defparam \fifo_data~218 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][14] (
	.clk(clk),
	.d(\fifo_data~218_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~201 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~201_combout ),
	.cout());
defparam \fifo_data~201 .lut_mask = 16'hEEEE;
defparam \fifo_data~201 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][14] (
	.clk(clk),
	.d(\fifo_data~201_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~184 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~184_combout ),
	.cout());
defparam \fifo_data~184 .lut_mask = 16'hEEEE;
defparam \fifo_data~184 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][14] (
	.clk(clk),
	.d(\fifo_data~184_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~167 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~167_combout ),
	.cout());
defparam \fifo_data~167 .lut_mask = 16'hEEEE;
defparam \fifo_data~167 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][14] (
	.clk(clk),
	.d(\fifo_data~167_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~150 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~150_combout ),
	.cout());
defparam \fifo_data~150 .lut_mask = 16'hEEEE;
defparam \fifo_data~150 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][14] (
	.clk(clk),
	.d(\fifo_data~150_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~133 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~133_combout ),
	.cout());
defparam \fifo_data~133 .lut_mask = 16'hEEEE;
defparam \fifo_data~133 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][14] (
	.clk(clk),
	.d(\fifo_data~133_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~116 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~116_combout ),
	.cout());
defparam \fifo_data~116 .lut_mask = 16'hEEEE;
defparam \fifo_data~116 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][14] (
	.clk(clk),
	.d(\fifo_data~116_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~99 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~99_combout ),
	.cout());
defparam \fifo_data~99 .lut_mask = 16'hEEEE;
defparam \fifo_data~99 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][14] (
	.clk(clk),
	.d(\fifo_data~99_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~82 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~82_combout ),
	.cout());
defparam \fifo_data~82 .lut_mask = 16'hEEEE;
defparam \fifo_data~82 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][14] (
	.clk(clk),
	.d(\fifo_data~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~65 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~65_combout ),
	.cout());
defparam \fifo_data~65 .lut_mask = 16'hEEEE;
defparam \fifo_data~65 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][14] (
	.clk(clk),
	.d(\fifo_data~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~48 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~48_combout ),
	.cout());
defparam \fifo_data~48 .lut_mask = 16'hEEEE;
defparam \fifo_data~48 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][14] (
	.clk(clk),
	.d(\fifo_data~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~31 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~31_combout ),
	.cout());
defparam \fifo_data~31 .lut_mask = 16'hEEEE;
defparam \fifo_data~31 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][14] (
	.clk(clk),
	.d(\fifo_data~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][14]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][14] .power_up = "low";

cycloneive_lcell_comb \fifo_data~14 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~14_combout ),
	.cout());
defparam \fifo_data~14 .lut_mask = 16'hEEEE;
defparam \fifo_data~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~270 (
	.dataa(reset_n),
	.datab(Mux1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~270_combout ),
	.cout());
defparam \fifo_data~270 .lut_mask = 16'hEEEE;
defparam \fifo_data~270 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\fifo_data~270_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~253 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~253_combout ),
	.cout());
defparam \fifo_data~253 .lut_mask = 16'hEEEE;
defparam \fifo_data~253 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][15] (
	.clk(clk),
	.d(\fifo_data~253_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~236 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~236_combout ),
	.cout());
defparam \fifo_data~236 .lut_mask = 16'hEEEE;
defparam \fifo_data~236 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][15] (
	.clk(clk),
	.d(\fifo_data~236_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~219 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~219_combout ),
	.cout());
defparam \fifo_data~219 .lut_mask = 16'hEEEE;
defparam \fifo_data~219 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][15] (
	.clk(clk),
	.d(\fifo_data~219_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~202 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~202_combout ),
	.cout());
defparam \fifo_data~202 .lut_mask = 16'hEEEE;
defparam \fifo_data~202 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][15] (
	.clk(clk),
	.d(\fifo_data~202_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~185 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~185_combout ),
	.cout());
defparam \fifo_data~185 .lut_mask = 16'hEEEE;
defparam \fifo_data~185 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][15] (
	.clk(clk),
	.d(\fifo_data~185_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~168 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~168_combout ),
	.cout());
defparam \fifo_data~168 .lut_mask = 16'hEEEE;
defparam \fifo_data~168 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][15] (
	.clk(clk),
	.d(\fifo_data~168_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~151 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~151_combout ),
	.cout());
defparam \fifo_data~151 .lut_mask = 16'hEEEE;
defparam \fifo_data~151 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][15] (
	.clk(clk),
	.d(\fifo_data~151_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~134 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~134_combout ),
	.cout());
defparam \fifo_data~134 .lut_mask = 16'hEEEE;
defparam \fifo_data~134 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][15] (
	.clk(clk),
	.d(\fifo_data~134_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~117 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~117_combout ),
	.cout());
defparam \fifo_data~117 .lut_mask = 16'hEEEE;
defparam \fifo_data~117 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][15] (
	.clk(clk),
	.d(\fifo_data~117_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~100 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~100_combout ),
	.cout());
defparam \fifo_data~100 .lut_mask = 16'hEEEE;
defparam \fifo_data~100 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][15] (
	.clk(clk),
	.d(\fifo_data~100_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~83 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~83_combout ),
	.cout());
defparam \fifo_data~83 .lut_mask = 16'hEEEE;
defparam \fifo_data~83 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][15] (
	.clk(clk),
	.d(\fifo_data~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~66 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~66_combout ),
	.cout());
defparam \fifo_data~66 .lut_mask = 16'hEEEE;
defparam \fifo_data~66 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][15] (
	.clk(clk),
	.d(\fifo_data~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~49 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~49_combout ),
	.cout());
defparam \fifo_data~49 .lut_mask = 16'hEEEE;
defparam \fifo_data~49 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][15] (
	.clk(clk),
	.d(\fifo_data~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~32 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~32_combout ),
	.cout());
defparam \fifo_data~32 .lut_mask = 16'hEEEE;
defparam \fifo_data~32 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][15] (
	.clk(clk),
	.d(\fifo_data~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][15]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][15] .power_up = "low";

cycloneive_lcell_comb \fifo_data~15 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~15_combout ),
	.cout());
defparam \fifo_data~15 .lut_mask = 16'hEEEE;
defparam \fifo_data~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_data~271 (
	.dataa(reset_n),
	.datab(Mux0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~271_combout ),
	.cout());
defparam \fifo_data~271 .lut_mask = 16'hEEEE;
defparam \fifo_data~271 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\fifo_data~271_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[0][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~254 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[0][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~254_combout ),
	.cout());
defparam \fifo_data~254 .lut_mask = 16'hEEEE;
defparam \fifo_data~254 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[1][16] (
	.clk(clk),
	.d(\fifo_data~254_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[1][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[1][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[1][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~237 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[1][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~237_combout ),
	.cout());
defparam \fifo_data~237 .lut_mask = 16'hEEEE;
defparam \fifo_data~237 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[2][16] (
	.clk(clk),
	.d(\fifo_data~237_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[2][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[2][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[2][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~220 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[2][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~220_combout ),
	.cout());
defparam \fifo_data~220 .lut_mask = 16'hEEEE;
defparam \fifo_data~220 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[3][16] (
	.clk(clk),
	.d(\fifo_data~220_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[3][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[3][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[3][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~203 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[3][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~203_combout ),
	.cout());
defparam \fifo_data~203 .lut_mask = 16'hEEEE;
defparam \fifo_data~203 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[4][16] (
	.clk(clk),
	.d(\fifo_data~203_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[4][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[4][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[4][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~186 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[4][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~186_combout ),
	.cout());
defparam \fifo_data~186 .lut_mask = 16'hEEEE;
defparam \fifo_data~186 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[5][16] (
	.clk(clk),
	.d(\fifo_data~186_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[5][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[5][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[5][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~169 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[5][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~169_combout ),
	.cout());
defparam \fifo_data~169 .lut_mask = 16'hEEEE;
defparam \fifo_data~169 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[6][16] (
	.clk(clk),
	.d(\fifo_data~169_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[6][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[6][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[6][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~152 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[6][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~152_combout ),
	.cout());
defparam \fifo_data~152 .lut_mask = 16'hEEEE;
defparam \fifo_data~152 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[7][16] (
	.clk(clk),
	.d(\fifo_data~152_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[7][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[7][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[7][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~135 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[7][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~135_combout ),
	.cout());
defparam \fifo_data~135 .lut_mask = 16'hEEEE;
defparam \fifo_data~135 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[8][16] (
	.clk(clk),
	.d(\fifo_data~135_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[8][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[8][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[8][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~118 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[8][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~118_combout ),
	.cout());
defparam \fifo_data~118 .lut_mask = 16'hEEEE;
defparam \fifo_data~118 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[9][16] (
	.clk(clk),
	.d(\fifo_data~118_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[9][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[9][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[9][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~101 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[9][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~101_combout ),
	.cout());
defparam \fifo_data~101 .lut_mask = 16'hEEEE;
defparam \fifo_data~101 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[10][16] (
	.clk(clk),
	.d(\fifo_data~101_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[10][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[10][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[10][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~84 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[10][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~84_combout ),
	.cout());
defparam \fifo_data~84 .lut_mask = 16'hEEEE;
defparam \fifo_data~84 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[11][16] (
	.clk(clk),
	.d(\fifo_data~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[11][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[11][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[11][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~67 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[11][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~67_combout ),
	.cout());
defparam \fifo_data~67 .lut_mask = 16'hEEEE;
defparam \fifo_data~67 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[12][16] (
	.clk(clk),
	.d(\fifo_data~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[12][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[12][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[12][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~50 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[12][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~50_combout ),
	.cout());
defparam \fifo_data~50 .lut_mask = 16'hEEEE;
defparam \fifo_data~50 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[13][16] (
	.clk(clk),
	.d(\fifo_data~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[13][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[13][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[13][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~33 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[13][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~33_combout ),
	.cout());
defparam \fifo_data~33 .lut_mask = 16'hEEEE;
defparam \fifo_data~33 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[14][16] (
	.clk(clk),
	.d(\fifo_data~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(register_fifofifo_data1414),
	.q(\register_fifo:fifo_data[14][16]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[14][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[14][16] .power_up = "low";

cycloneive_lcell_comb \fifo_data~16 (
	.dataa(reset_n),
	.datab(\register_fifo:fifo_data[14][16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_data~16_combout ),
	.cout());
defparam \fifo_data~16 .lut_mask = 16'hEEEE;
defparam \fifo_data~16 .sum_lutc_input = "datac";

endmodule

module CIC_auk_dspip_downsample (
	sample_state_0,
	count_0,
	count_3,
	count_4,
	count_2,
	count_5,
	count_6,
	count_7,
	count_8,
	count_9,
	count_1,
	stall_reg,
	ena_sample,
	Equal0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	count_0;
output 	count_3;
output 	count_4;
output 	count_2;
output 	count_5;
output 	count_6;
output 	count_7;
output 	count_8;
output 	count_9;
output 	count_1;
input 	stall_reg;
input 	ena_sample;
output 	Equal0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_counter_module_1 counter_fs_inst(
	.sample_state_0(sample_state_0),
	.count_0(count_0),
	.count_3(count_3),
	.count_4(count_4),
	.count_2(count_2),
	.count_5(count_5),
	.count_6(count_6),
	.count_7(count_7),
	.count_8(count_8),
	.count_9(count_9),
	.count_1(count_1),
	.stall_reg(stall_reg),
	.ena_sample(ena_sample),
	.Equal0(Equal0),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_counter_module_1 (
	sample_state_0,
	count_0,
	count_3,
	count_4,
	count_2,
	count_5,
	count_6,
	count_7,
	count_8,
	count_9,
	count_1,
	stall_reg,
	ena_sample,
	Equal0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	count_0;
output 	count_3;
output 	count_4;
output 	count_2;
output 	count_5;
output 	count_6;
output 	count_7;
output 	count_8;
output 	count_9;
output 	count_1;
input 	stall_reg;
input 	ena_sample;
output 	Equal0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \count[0]~10_combout ;
wire \Equal0~1_combout ;
wire \count[5]~12_combout ;
wire \count[5]~13_combout ;
wire \count[0]~11 ;
wire \count[1]~15 ;
wire \count[2]~17 ;
wire \count[3]~18_combout ;
wire \count[3]~19 ;
wire \count[4]~20_combout ;
wire \count[2]~16_combout ;
wire \count[4]~21 ;
wire \count[5]~22_combout ;
wire \count[5]~23 ;
wire \count[6]~24_combout ;
wire \count[6]~25 ;
wire \count[7]~26_combout ;
wire \count[7]~27 ;
wire \count[8]~28_combout ;
wire \count[8]~29 ;
wire \count[9]~30_combout ;
wire \count[1]~14_combout ;


dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_3),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_4),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_2),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_5),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_6),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[7] (
	.clk(clk),
	.d(\count[7]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_7),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

dffeas \count[8] (
	.clk(clk),
	.d(\count[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_8),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

dffeas \count[9] (
	.clk(clk),
	.d(\count[9]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_9),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[5]~12_combout ),
	.sload(gnd),
	.ena(\count[5]~13_combout ),
	.q(count_1),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(count_5),
	.datab(count_6),
	.datac(count_7),
	.datad(count_8),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFFFE;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[0]~10 (
	.dataa(count_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~10_combout ),
	.cout(\count[0]~11 ));
defparam \count[0]~10 .lut_mask = 16'h55AA;
defparam \count[0]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(count_1),
	.datab(count_0),
	.datac(ena_sample),
	.datad(count_2),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h7FFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[5]~12 (
	.dataa(reset_n),
	.datab(\Equal0~1_combout ),
	.datac(count_9),
	.datad(Equal0),
	.cin(gnd),
	.combout(\count[5]~12_combout ),
	.cout());
defparam \count[5]~12 .lut_mask = 16'hFFF7;
defparam \count[5]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[5]~13 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(sample_state_0),
	.cin(gnd),
	.combout(\count[5]~13_combout ),
	.cout());
defparam \count[5]~13 .lut_mask = 16'hFF77;
defparam \count[5]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[1]~14 (
	.dataa(count_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~11 ),
	.combout(\count[1]~14_combout ),
	.cout(\count[1]~15 ));
defparam \count[1]~14 .lut_mask = 16'h5A5F;
defparam \count[1]~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[2]~16 (
	.dataa(count_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~15 ),
	.combout(\count[2]~16_combout ),
	.cout(\count[2]~17 ));
defparam \count[2]~16 .lut_mask = 16'h5AAF;
defparam \count[2]~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[3]~18 (
	.dataa(count_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~17 ),
	.combout(\count[3]~18_combout ),
	.cout(\count[3]~19 ));
defparam \count[3]~18 .lut_mask = 16'h5A5F;
defparam \count[3]~18 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[4]~20 (
	.dataa(count_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~19 ),
	.combout(\count[4]~20_combout ),
	.cout(\count[4]~21 ));
defparam \count[4]~20 .lut_mask = 16'h5AAF;
defparam \count[4]~20 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[5]~22 (
	.dataa(count_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~21 ),
	.combout(\count[5]~22_combout ),
	.cout(\count[5]~23 ));
defparam \count[5]~22 .lut_mask = 16'h5A5F;
defparam \count[5]~22 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[6]~24 (
	.dataa(count_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[5]~23 ),
	.combout(\count[6]~24_combout ),
	.cout(\count[6]~25 ));
defparam \count[6]~24 .lut_mask = 16'h5AAF;
defparam \count[6]~24 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[7]~26 (
	.dataa(count_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[6]~25 ),
	.combout(\count[7]~26_combout ),
	.cout(\count[7]~27 ));
defparam \count[7]~26 .lut_mask = 16'h5A5F;
defparam \count[7]~26 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[8]~28 (
	.dataa(count_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[7]~27 ),
	.combout(\count[8]~28_combout ),
	.cout(\count[8]~29 ));
defparam \count[8]~28 .lut_mask = 16'h5AAF;
defparam \count[8]~28 .sum_lutc_input = "cin";

cycloneive_lcell_comb \count[9]~30 (
	.dataa(count_9),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[8]~29 ),
	.combout(\count[9]~30_combout ),
	.cout());
defparam \count[9]~30 .lut_mask = 16'h5A5A;
defparam \count[9]~30 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	stall_reg,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_10;
input 	q_b_9;
input 	q_b_8;
input 	q_b_7;
input 	q_b_6;
input 	q_b_5;
input 	q_b_4;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	stall_reg;
output 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_1 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_10(q_b_10),
	.q_b_9(q_b_9),
	.q_b_8(q_b_8),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.stall_reg(stall_reg),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_1 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	stall_reg,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_10;
input 	q_b_9;
input 	q_b_8;
input 	q_b_7;
input 	q_b_6;
input 	q_b_5;
input 	q_b_4;
input 	q_b_11;
input 	q_b_12;
input 	q_b_13;
input 	q_b_14;
input 	q_b_15;
input 	stall_reg;
output 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~2_combout ;
wire \register_fifo:fifo_data[0][13]~3 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(register_fifofifo_data0131),
	.cout());
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h7777;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~2 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~2_combout ),
	.cout(\register_fifo:fifo_data[0][13]~3 ));
defparam \register_fifo:fifo_data[0][13]~2 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~3 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_15),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_1 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_170,
	q_b_169,
	q_b_168,
	q_b_167,
	q_b_166,
	q_b_165,
	q_b_164,
	q_b_171,
	q_b_172,
	q_b_173,
	q_b_174,
	q_b_175,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_170;
input 	q_b_169;
input 	q_b_168;
input 	q_b_167;
input 	q_b_166;
input 	q_b_165;
input 	q_b_164;
input 	q_b_171;
input 	q_b_172;
input 	q_b_173;
input 	q_b_174;
input 	q_b_175;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_2 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_170(q_b_170),
	.q_b_169(q_b_169),
	.q_b_168(q_b_168),
	.q_b_167(q_b_167),
	.q_b_166(q_b_166),
	.q_b_165(q_b_165),
	.q_b_164(q_b_164),
	.q_b_171(q_b_171),
	.q_b_172(q_b_172),
	.q_b_173(q_b_173),
	.q_b_174(q_b_174),
	.q_b_175(q_b_175),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_2 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_170,
	q_b_169,
	q_b_168,
	q_b_167,
	q_b_166,
	q_b_165,
	q_b_164,
	q_b_171,
	q_b_172,
	q_b_173,
	q_b_174,
	q_b_175,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_170;
input 	q_b_169;
input 	q_b_168;
input 	q_b_167;
input 	q_b_166;
input 	q_b_165;
input 	q_b_164;
input 	q_b_171;
input 	q_b_172;
input 	q_b_173;
input 	q_b_174;
input 	q_b_175;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_164),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_165),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_166),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_167),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_168),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_169),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_170),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_172),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_173),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_174),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_175),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_175),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_2 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_186,
	q_b_185,
	q_b_184,
	q_b_183,
	q_b_182,
	q_b_181,
	q_b_180,
	q_b_187,
	q_b_188,
	q_b_189,
	q_b_190,
	q_b_191,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_186;
input 	q_b_185;
input 	q_b_184;
input 	q_b_183;
input 	q_b_182;
input 	q_b_181;
input 	q_b_180;
input 	q_b_187;
input 	q_b_188;
input 	q_b_189;
input 	q_b_190;
input 	q_b_191;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_3 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_186(q_b_186),
	.q_b_185(q_b_185),
	.q_b_184(q_b_184),
	.q_b_183(q_b_183),
	.q_b_182(q_b_182),
	.q_b_181(q_b_181),
	.q_b_180(q_b_180),
	.q_b_187(q_b_187),
	.q_b_188(q_b_188),
	.q_b_189(q_b_189),
	.q_b_190(q_b_190),
	.q_b_191(q_b_191),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_3 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_186,
	q_b_185,
	q_b_184,
	q_b_183,
	q_b_182,
	q_b_181,
	q_b_180,
	q_b_187,
	q_b_188,
	q_b_189,
	q_b_190,
	q_b_191,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_186;
input 	q_b_185;
input 	q_b_184;
input 	q_b_183;
input 	q_b_182;
input 	q_b_181;
input 	q_b_180;
input 	q_b_187;
input 	q_b_188;
input 	q_b_189;
input 	q_b_190;
input 	q_b_191;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_180),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_181),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_182),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_183),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_184),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_185),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_186),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_187),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_188),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_189),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_190),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_191),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_191),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_3 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_202,
	q_b_201,
	q_b_200,
	q_b_199,
	q_b_198,
	q_b_197,
	q_b_196,
	q_b_203,
	q_b_204,
	q_b_205,
	q_b_206,
	q_b_207,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_202;
input 	q_b_201;
input 	q_b_200;
input 	q_b_199;
input 	q_b_198;
input 	q_b_197;
input 	q_b_196;
input 	q_b_203;
input 	q_b_204;
input 	q_b_205;
input 	q_b_206;
input 	q_b_207;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_4 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_202(q_b_202),
	.q_b_201(q_b_201),
	.q_b_200(q_b_200),
	.q_b_199(q_b_199),
	.q_b_198(q_b_198),
	.q_b_197(q_b_197),
	.q_b_196(q_b_196),
	.q_b_203(q_b_203),
	.q_b_204(q_b_204),
	.q_b_205(q_b_205),
	.q_b_206(q_b_206),
	.q_b_207(q_b_207),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_4 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_202,
	q_b_201,
	q_b_200,
	q_b_199,
	q_b_198,
	q_b_197,
	q_b_196,
	q_b_203,
	q_b_204,
	q_b_205,
	q_b_206,
	q_b_207,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_202;
input 	q_b_201;
input 	q_b_200;
input 	q_b_199;
input 	q_b_198;
input 	q_b_197;
input 	q_b_196;
input 	q_b_203;
input 	q_b_204;
input 	q_b_205;
input 	q_b_206;
input 	q_b_207;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_196),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_197),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_198),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_199),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_200),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_201),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_202),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_203),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_204),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_205),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_206),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_207),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_207),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_4 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_218,
	q_b_217,
	q_b_216,
	q_b_215,
	q_b_214,
	q_b_213,
	q_b_212,
	q_b_219,
	q_b_220,
	q_b_221,
	q_b_222,
	q_b_223,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_218;
input 	q_b_217;
input 	q_b_216;
input 	q_b_215;
input 	q_b_214;
input 	q_b_213;
input 	q_b_212;
input 	q_b_219;
input 	q_b_220;
input 	q_b_221;
input 	q_b_222;
input 	q_b_223;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_5 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_218(q_b_218),
	.q_b_217(q_b_217),
	.q_b_216(q_b_216),
	.q_b_215(q_b_215),
	.q_b_214(q_b_214),
	.q_b_213(q_b_213),
	.q_b_212(q_b_212),
	.q_b_219(q_b_219),
	.q_b_220(q_b_220),
	.q_b_221(q_b_221),
	.q_b_222(q_b_222),
	.q_b_223(q_b_223),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_5 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_218,
	q_b_217,
	q_b_216,
	q_b_215,
	q_b_214,
	q_b_213,
	q_b_212,
	q_b_219,
	q_b_220,
	q_b_221,
	q_b_222,
	q_b_223,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_218;
input 	q_b_217;
input 	q_b_216;
input 	q_b_215;
input 	q_b_214;
input 	q_b_213;
input 	q_b_212;
input 	q_b_219;
input 	q_b_220;
input 	q_b_221;
input 	q_b_222;
input 	q_b_223;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_212),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_213),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_214),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_215),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_216),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_217),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_218),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_219),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_220),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_221),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_222),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_223),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_223),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_5 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_234,
	q_b_233,
	q_b_232,
	q_b_231,
	q_b_230,
	q_b_229,
	q_b_228,
	q_b_235,
	q_b_236,
	q_b_237,
	q_b_238,
	q_b_239,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_234;
input 	q_b_233;
input 	q_b_232;
input 	q_b_231;
input 	q_b_230;
input 	q_b_229;
input 	q_b_228;
input 	q_b_235;
input 	q_b_236;
input 	q_b_237;
input 	q_b_238;
input 	q_b_239;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_6 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_234(q_b_234),
	.q_b_233(q_b_233),
	.q_b_232(q_b_232),
	.q_b_231(q_b_231),
	.q_b_230(q_b_230),
	.q_b_229(q_b_229),
	.q_b_228(q_b_228),
	.q_b_235(q_b_235),
	.q_b_236(q_b_236),
	.q_b_237(q_b_237),
	.q_b_238(q_b_238),
	.q_b_239(q_b_239),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_6 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_234,
	q_b_233,
	q_b_232,
	q_b_231,
	q_b_230,
	q_b_229,
	q_b_228,
	q_b_235,
	q_b_236,
	q_b_237,
	q_b_238,
	q_b_239,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_234;
input 	q_b_233;
input 	q_b_232;
input 	q_b_231;
input 	q_b_230;
input 	q_b_229;
input 	q_b_228;
input 	q_b_235;
input 	q_b_236;
input 	q_b_237;
input 	q_b_238;
input 	q_b_239;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_228),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_229),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_230),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_231),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_232),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_233),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_234),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_235),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_236),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_237),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_238),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_239),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_239),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_6 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_250,
	q_b_249,
	q_b_248,
	q_b_247,
	q_b_246,
	q_b_245,
	q_b_244,
	q_b_251,
	q_b_252,
	q_b_253,
	q_b_254,
	q_b_255,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_250;
input 	q_b_249;
input 	q_b_248;
input 	q_b_247;
input 	q_b_246;
input 	q_b_245;
input 	q_b_244;
input 	q_b_251;
input 	q_b_252;
input 	q_b_253;
input 	q_b_254;
input 	q_b_255;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_7 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_250(q_b_250),
	.q_b_249(q_b_249),
	.q_b_248(q_b_248),
	.q_b_247(q_b_247),
	.q_b_246(q_b_246),
	.q_b_245(q_b_245),
	.q_b_244(q_b_244),
	.q_b_251(q_b_251),
	.q_b_252(q_b_252),
	.q_b_253(q_b_253),
	.q_b_254(q_b_254),
	.q_b_255(q_b_255),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_7 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_250,
	q_b_249,
	q_b_248,
	q_b_247,
	q_b_246,
	q_b_245,
	q_b_244,
	q_b_251,
	q_b_252,
	q_b_253,
	q_b_254,
	q_b_255,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_250;
input 	q_b_249;
input 	q_b_248;
input 	q_b_247;
input 	q_b_246;
input 	q_b_245;
input 	q_b_244;
input 	q_b_251;
input 	q_b_252;
input 	q_b_253;
input 	q_b_254;
input 	q_b_255;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_244),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_245),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_246),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_247),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_248),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_249),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_250),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_251),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_252),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_253),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_254),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_255),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_255),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_7 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_26;
input 	q_b_25;
input 	q_b_24;
input 	q_b_23;
input 	q_b_22;
input 	q_b_21;
input 	q_b_20;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_8 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_26(q_b_26),
	.q_b_25(q_b_25),
	.q_b_24(q_b_24),
	.q_b_23(q_b_23),
	.q_b_22(q_b_22),
	.q_b_21(q_b_21),
	.q_b_20(q_b_20),
	.q_b_27(q_b_27),
	.q_b_28(q_b_28),
	.q_b_29(q_b_29),
	.q_b_30(q_b_30),
	.q_b_31(q_b_31),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_8 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_26,
	q_b_25,
	q_b_24,
	q_b_23,
	q_b_22,
	q_b_21,
	q_b_20,
	q_b_27,
	q_b_28,
	q_b_29,
	q_b_30,
	q_b_31,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_26;
input 	q_b_25;
input 	q_b_24;
input 	q_b_23;
input 	q_b_22;
input 	q_b_21;
input 	q_b_20;
input 	q_b_27;
input 	q_b_28;
input 	q_b_29;
input 	q_b_30;
input 	q_b_31;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_20),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_28),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_31),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_8 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_42,
	q_b_41,
	q_b_40,
	q_b_39,
	q_b_38,
	q_b_37,
	q_b_36,
	q_b_43,
	q_b_44,
	q_b_45,
	q_b_46,
	q_b_47,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_42;
input 	q_b_41;
input 	q_b_40;
input 	q_b_39;
input 	q_b_38;
input 	q_b_37;
input 	q_b_36;
input 	q_b_43;
input 	q_b_44;
input 	q_b_45;
input 	q_b_46;
input 	q_b_47;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_9 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_42(q_b_42),
	.q_b_41(q_b_41),
	.q_b_40(q_b_40),
	.q_b_39(q_b_39),
	.q_b_38(q_b_38),
	.q_b_37(q_b_37),
	.q_b_36(q_b_36),
	.q_b_43(q_b_43),
	.q_b_44(q_b_44),
	.q_b_45(q_b_45),
	.q_b_46(q_b_46),
	.q_b_47(q_b_47),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_9 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_42,
	q_b_41,
	q_b_40,
	q_b_39,
	q_b_38,
	q_b_37,
	q_b_36,
	q_b_43,
	q_b_44,
	q_b_45,
	q_b_46,
	q_b_47,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_42;
input 	q_b_41;
input 	q_b_40;
input 	q_b_39;
input 	q_b_38;
input 	q_b_37;
input 	q_b_36;
input 	q_b_43;
input 	q_b_44;
input 	q_b_45;
input 	q_b_46;
input 	q_b_47;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_36),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_37),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_38),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_39),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_40),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_42),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_43),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_44),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_45),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_46),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_47),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_47),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_9 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_58,
	q_b_57,
	q_b_56,
	q_b_55,
	q_b_54,
	q_b_53,
	q_b_52,
	q_b_59,
	q_b_60,
	q_b_61,
	q_b_62,
	q_b_63,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_58;
input 	q_b_57;
input 	q_b_56;
input 	q_b_55;
input 	q_b_54;
input 	q_b_53;
input 	q_b_52;
input 	q_b_59;
input 	q_b_60;
input 	q_b_61;
input 	q_b_62;
input 	q_b_63;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_10 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_58(q_b_58),
	.q_b_57(q_b_57),
	.q_b_56(q_b_56),
	.q_b_55(q_b_55),
	.q_b_54(q_b_54),
	.q_b_53(q_b_53),
	.q_b_52(q_b_52),
	.q_b_59(q_b_59),
	.q_b_60(q_b_60),
	.q_b_61(q_b_61),
	.q_b_62(q_b_62),
	.q_b_63(q_b_63),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_10 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_58,
	q_b_57,
	q_b_56,
	q_b_55,
	q_b_54,
	q_b_53,
	q_b_52,
	q_b_59,
	q_b_60,
	q_b_61,
	q_b_62,
	q_b_63,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_58;
input 	q_b_57;
input 	q_b_56;
input 	q_b_55;
input 	q_b_54;
input 	q_b_53;
input 	q_b_52;
input 	q_b_59;
input 	q_b_60;
input 	q_b_61;
input 	q_b_62;
input 	q_b_63;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_52),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_53),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_54),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_55),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_56),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_57),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_58),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_59),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_60),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_61),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_62),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_63),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_63),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_10 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_74,
	q_b_73,
	q_b_72,
	q_b_71,
	q_b_70,
	q_b_69,
	q_b_68,
	q_b_75,
	q_b_76,
	q_b_77,
	q_b_78,
	q_b_79,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_74;
input 	q_b_73;
input 	q_b_72;
input 	q_b_71;
input 	q_b_70;
input 	q_b_69;
input 	q_b_68;
input 	q_b_75;
input 	q_b_76;
input 	q_b_77;
input 	q_b_78;
input 	q_b_79;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_11 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_74(q_b_74),
	.q_b_73(q_b_73),
	.q_b_72(q_b_72),
	.q_b_71(q_b_71),
	.q_b_70(q_b_70),
	.q_b_69(q_b_69),
	.q_b_68(q_b_68),
	.q_b_75(q_b_75),
	.q_b_76(q_b_76),
	.q_b_77(q_b_77),
	.q_b_78(q_b_78),
	.q_b_79(q_b_79),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_11 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_74,
	q_b_73,
	q_b_72,
	q_b_71,
	q_b_70,
	q_b_69,
	q_b_68,
	q_b_75,
	q_b_76,
	q_b_77,
	q_b_78,
	q_b_79,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_74;
input 	q_b_73;
input 	q_b_72;
input 	q_b_71;
input 	q_b_70;
input 	q_b_69;
input 	q_b_68;
input 	q_b_75;
input 	q_b_76;
input 	q_b_77;
input 	q_b_78;
input 	q_b_79;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_68),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_69),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_70),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_71),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_72),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_73),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_74),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_75),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_76),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_77),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_78),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_79),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_79),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_11 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_90,
	q_b_89,
	q_b_88,
	q_b_87,
	q_b_86,
	q_b_85,
	q_b_84,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_94,
	q_b_95,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_90;
input 	q_b_89;
input 	q_b_88;
input 	q_b_87;
input 	q_b_86;
input 	q_b_85;
input 	q_b_84;
input 	q_b_91;
input 	q_b_92;
input 	q_b_93;
input 	q_b_94;
input 	q_b_95;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_12 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_90(q_b_90),
	.q_b_89(q_b_89),
	.q_b_88(q_b_88),
	.q_b_87(q_b_87),
	.q_b_86(q_b_86),
	.q_b_85(q_b_85),
	.q_b_84(q_b_84),
	.q_b_91(q_b_91),
	.q_b_92(q_b_92),
	.q_b_93(q_b_93),
	.q_b_94(q_b_94),
	.q_b_95(q_b_95),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_12 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_90,
	q_b_89,
	q_b_88,
	q_b_87,
	q_b_86,
	q_b_85,
	q_b_84,
	q_b_91,
	q_b_92,
	q_b_93,
	q_b_94,
	q_b_95,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_90;
input 	q_b_89;
input 	q_b_88;
input 	q_b_87;
input 	q_b_86;
input 	q_b_85;
input 	q_b_84;
input 	q_b_91;
input 	q_b_92;
input 	q_b_93;
input 	q_b_94;
input 	q_b_95;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_84),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_85),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_86),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_87),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_88),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_89),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_90),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_91),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_92),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_93),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_94),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_95),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_95),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_12 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_106,
	q_b_105,
	q_b_104,
	q_b_103,
	q_b_102,
	q_b_101,
	q_b_100,
	q_b_107,
	q_b_108,
	q_b_109,
	q_b_110,
	q_b_111,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_106;
input 	q_b_105;
input 	q_b_104;
input 	q_b_103;
input 	q_b_102;
input 	q_b_101;
input 	q_b_100;
input 	q_b_107;
input 	q_b_108;
input 	q_b_109;
input 	q_b_110;
input 	q_b_111;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_13 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_106(q_b_106),
	.q_b_105(q_b_105),
	.q_b_104(q_b_104),
	.q_b_103(q_b_103),
	.q_b_102(q_b_102),
	.q_b_101(q_b_101),
	.q_b_100(q_b_100),
	.q_b_107(q_b_107),
	.q_b_108(q_b_108),
	.q_b_109(q_b_109),
	.q_b_110(q_b_110),
	.q_b_111(q_b_111),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_13 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_106,
	q_b_105,
	q_b_104,
	q_b_103,
	q_b_102,
	q_b_101,
	q_b_100,
	q_b_107,
	q_b_108,
	q_b_109,
	q_b_110,
	q_b_111,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_106;
input 	q_b_105;
input 	q_b_104;
input 	q_b_103;
input 	q_b_102;
input 	q_b_101;
input 	q_b_100;
input 	q_b_107;
input 	q_b_108;
input 	q_b_109;
input 	q_b_110;
input 	q_b_111;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_100),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_102),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_103),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_104),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_105),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_106),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_107),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_108),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_109),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_110),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_111),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_13 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_122,
	q_b_121,
	q_b_120,
	q_b_119,
	q_b_118,
	q_b_117,
	q_b_116,
	q_b_123,
	q_b_124,
	q_b_125,
	q_b_126,
	q_b_127,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_122;
input 	q_b_121;
input 	q_b_120;
input 	q_b_119;
input 	q_b_118;
input 	q_b_117;
input 	q_b_116;
input 	q_b_123;
input 	q_b_124;
input 	q_b_125;
input 	q_b_126;
input 	q_b_127;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_14 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_122(q_b_122),
	.q_b_121(q_b_121),
	.q_b_120(q_b_120),
	.q_b_119(q_b_119),
	.q_b_118(q_b_118),
	.q_b_117(q_b_117),
	.q_b_116(q_b_116),
	.q_b_123(q_b_123),
	.q_b_124(q_b_124),
	.q_b_125(q_b_125),
	.q_b_126(q_b_126),
	.q_b_127(q_b_127),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_14 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_122,
	q_b_121,
	q_b_120,
	q_b_119,
	q_b_118,
	q_b_117,
	q_b_116,
	q_b_123,
	q_b_124,
	q_b_125,
	q_b_126,
	q_b_127,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_122;
input 	q_b_121;
input 	q_b_120;
input 	q_b_119;
input 	q_b_118;
input 	q_b_117;
input 	q_b_116;
input 	q_b_123;
input 	q_b_124;
input 	q_b_125;
input 	q_b_126;
input 	q_b_127;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_116),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_117),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_118),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_119),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_120),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_122),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_123),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_124),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_125),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_126),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_127),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_127),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_14 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_138,
	q_b_137,
	q_b_136,
	q_b_135,
	q_b_134,
	q_b_133,
	q_b_132,
	q_b_139,
	q_b_140,
	q_b_141,
	q_b_142,
	q_b_143,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_138;
input 	q_b_137;
input 	q_b_136;
input 	q_b_135;
input 	q_b_134;
input 	q_b_133;
input 	q_b_132;
input 	q_b_139;
input 	q_b_140;
input 	q_b_141;
input 	q_b_142;
input 	q_b_143;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_15 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_138(q_b_138),
	.q_b_137(q_b_137),
	.q_b_136(q_b_136),
	.q_b_135(q_b_135),
	.q_b_134(q_b_134),
	.q_b_133(q_b_133),
	.q_b_132(q_b_132),
	.q_b_139(q_b_139),
	.q_b_140(q_b_140),
	.q_b_141(q_b_141),
	.q_b_142(q_b_142),
	.q_b_143(q_b_143),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_15 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_138,
	q_b_137,
	q_b_136,
	q_b_135,
	q_b_134,
	q_b_133,
	q_b_132,
	q_b_139,
	q_b_140,
	q_b_141,
	q_b_142,
	q_b_143,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_138;
input 	q_b_137;
input 	q_b_136;
input 	q_b_135;
input 	q_b_134;
input 	q_b_133;
input 	q_b_132;
input 	q_b_139;
input 	q_b_140;
input 	q_b_141;
input 	q_b_142;
input 	q_b_143;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_132),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_133),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_134),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_135),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_136),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_137),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_138),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_139),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_140),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_142),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_143),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_143),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_integrator_15 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_154,
	q_b_153,
	q_b_152,
	q_b_151,
	q_b_150,
	q_b_149,
	q_b_148,
	q_b_155,
	q_b_156,
	q_b_157,
	q_b_158,
	q_b_159,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_154;
input 	q_b_153;
input 	q_b_152;
input 	q_b_151;
input 	q_b_150;
input 	q_b_149;
input 	q_b_148;
input 	q_b_155;
input 	q_b_156;
input 	q_b_157;
input 	q_b_158;
input 	q_b_159;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_auk_dspip_delay_16 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data020(register_fifofifo_data020),
	.register_fifofifo_data021(register_fifofifo_data021),
	.q_b_154(q_b_154),
	.q_b_153(q_b_153),
	.q_b_152(q_b_152),
	.q_b_151(q_b_151),
	.q_b_150(q_b_150),
	.q_b_149(q_b_149),
	.q_b_148(q_b_148),
	.q_b_155(q_b_155),
	.q_b_156(q_b_156),
	.q_b_157(q_b_157),
	.q_b_158(q_b_158),
	.q_b_159(q_b_159),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module CIC_auk_dspip_delay_16 (
	register_fifofifo_data06,
	register_fifofifo_data05,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data019,
	register_fifofifo_data020,
	register_fifofifo_data021,
	q_b_154,
	q_b_153,
	q_b_152,
	q_b_151,
	q_b_150,
	q_b_149,
	q_b_148,
	q_b_155,
	q_b_156,
	q_b_157,
	q_b_158,
	q_b_159,
	register_fifofifo_data0131,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data06;
output 	register_fifofifo_data05;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
output 	register_fifofifo_data019;
output 	register_fifofifo_data020;
output 	register_fifofifo_data021;
input 	q_b_154;
input 	q_b_153;
input 	q_b_152;
input 	q_b_151;
input 	q_b_150;
input 	q_b_149;
input 	q_b_148;
input 	q_b_155;
input 	q_b_156;
input 	q_b_157;
input 	q_b_158;
input 	q_b_159;
input 	register_fifofifo_data0131;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~q ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~q ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~q ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~q ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~q ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;
wire \register_fifo:fifo_data[0][18]~2 ;
wire \register_fifo:fifo_data[0][19]~1_combout ;
wire \register_fifo:fifo_data[0][19]~2 ;
wire \register_fifo:fifo_data[0][20]~1_combout ;
wire \register_fifo:fifo_data[0][20]~2 ;
wire \register_fifo:fifo_data[0][21]~1_combout ;


dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

dffeas \register_fifo:fifo_data[0][19] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][19]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data019),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][19] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][19] .power_up = "low";

dffeas \register_fifo:fifo_data[0][20] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][20]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data020),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][20] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][20] .power_up = "low";

dffeas \register_fifo:fifo_data[0][21] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][21]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(register_fifofifo_data021),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][21] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][21] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(\register_fifo:fifo_data[0][0]~q ),
	.datab(q_b_148),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(\register_fifo:fifo_data[0][1]~q ),
	.datab(q_b_149),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(\register_fifo:fifo_data[0][2]~q ),
	.datab(q_b_150),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(\register_fifo:fifo_data[0][3]~q ),
	.datab(q_b_151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][3]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(\register_fifo:fifo_data[0][4]~q ),
	.datab(q_b_152),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(register_fifofifo_data0131),
	.q(\register_fifo:fifo_data[0][4]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

cycloneive_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_153),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_154),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_155),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_156),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_157),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_158),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout(\register_fifo:fifo_data[0][18]~2 ));
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][19]~1 (
	.dataa(register_fifofifo_data019),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]~2 ),
	.combout(\register_fifo:fifo_data[0][19]~1_combout ),
	.cout(\register_fifo:fifo_data[0][19]~2 ));
defparam \register_fifo:fifo_data[0][19]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][19]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][20]~1 (
	.dataa(register_fifofifo_data020),
	.datab(q_b_159),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][19]~2 ),
	.combout(\register_fifo:fifo_data[0][20]~1_combout ),
	.cout(\register_fifo:fifo_data[0][20]~2 ));
defparam \register_fifo:fifo_data[0][20]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][20]~1 .sum_lutc_input = "cin";

cycloneive_lcell_comb \register_fifo:fifo_data[0][21]~1 (
	.dataa(register_fifofifo_data021),
	.datab(q_b_159),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][20]~2 ),
	.combout(\register_fifo:fifo_data[0][21]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][21]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][21]~1 .sum_lutc_input = "cin";

endmodule

module CIC_counter_module_33 (
	ena_sample,
	stall_reg,
	count_1,
	count_0,
	count_2,
	count_3,
	Equal6,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	ena_sample;
input 	stall_reg;
output 	count_1;
output 	count_0;
output 	count_2;
output 	count_3;
input 	Equal6;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \count~6_combout ;
wire \count[0]~2_combout ;
wire \count~3_combout ;
wire \Add0~0_combout ;
wire \count~4_combout ;
wire \Add0~1_combout ;
wire \count~5_combout ;


dffeas \count[1] (
	.clk(clk),
	.d(\count~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_1),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

dffeas \count[0] (
	.clk(clk),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_2),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_3),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

cycloneive_lcell_comb \count~6 (
	.dataa(count_1),
	.datab(count_0),
	.datac(reset_n),
	.datad(Equal6),
	.cin(gnd),
	.combout(\count~6_combout ),
	.cout());
defparam \count~6 .lut_mask = 16'hF6FF;
defparam \count~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count[0]~2 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(ena_sample),
	.cin(gnd),
	.combout(\count[0]~2_combout ),
	.cout());
defparam \count[0]~2 .lut_mask = 16'hFF77;
defparam \count[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count~3 (
	.dataa(count_0),
	.datab(Equal6),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
defparam \count~3 .lut_mask = 16'hFF77;
defparam \count~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(count_2),
	.datac(count_1),
	.datad(count_0),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'hC33C;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count~4 (
	.dataa(reset_n),
	.datab(\Add0~0_combout ),
	.datac(gnd),
	.datad(Equal6),
	.cin(gnd),
	.combout(\count~4_combout ),
	.cout());
defparam \count~4 .lut_mask = 16'hEEFF;
defparam \count~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~1 (
	.dataa(count_3),
	.datab(count_2),
	.datac(count_1),
	.datad(count_0),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'h6996;
defparam \Add0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \count~5 (
	.dataa(reset_n),
	.datab(\Add0~1_combout ),
	.datac(gnd),
	.datad(Equal6),
	.cin(gnd),
	.combout(\count~5_combout ),
	.cout());
defparam \count~5 .lut_mask = 16'hEEFF;
defparam \count~5 .sum_lutc_input = "datac";

endmodule

module CIC_auk_dspip_avalon_streaming_controller (
	dffe_nae,
	dffe_af,
	sink_ready_ctrl,
	stall_reg1,
	usedw_process,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	dffe_nae;
input 	dffe_af;
output 	sink_ready_ctrl;
output 	stall_reg1;
output 	usedw_process;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ready_FIFO|fifo_array[5][0]~q ;
wire \ready_FIFO|fifo_array[4][0]~q ;
wire \ready_FIFO|rd_addr_ptr[2]~q ;
wire \ready_FIFO|rd_addr_ptr[0]~q ;
wire \ready_FIFO|rd_addr_ptr[1]~q ;
wire \ready_FIFO|Equal2~0_combout ;
wire \ready_FIFO|Mux0~1_combout ;
wire \sink_ready_ctrl~0_combout ;
wire \sink_ready_ctrl~1_combout ;
wire \stall_reg~0_combout ;


CIC_auk_dspip_avalon_streaming_small_fifo ready_FIFO(
	.dffe_nae(dffe_nae),
	.fifo_array_0_5(\ready_FIFO|fifo_array[5][0]~q ),
	.fifo_array_0_4(\ready_FIFO|fifo_array[4][0]~q ),
	.rd_addr_ptr_2(\ready_FIFO|rd_addr_ptr[2]~q ),
	.dffe_af(dffe_af),
	.rd_addr_ptr_0(\ready_FIFO|rd_addr_ptr[0]~q ),
	.rd_addr_ptr_1(\ready_FIFO|rd_addr_ptr[1]~q ),
	.Equal2(\ready_FIFO|Equal2~0_combout ),
	.Mux0(\ready_FIFO|Mux0~1_combout ),
	.stall_reg(stall_reg1),
	.usedw_process(usedw_process),
	.clock(clk),
	.reset_n(reset_n));

cycloneive_lcell_comb \sink_ready_ctrl~2 (
	.dataa(\sink_ready_ctrl~1_combout ),
	.datab(\ready_FIFO|Equal2~0_combout ),
	.datac(\ready_FIFO|Mux0~1_combout ),
	.datad(\ready_FIFO|rd_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(sink_ready_ctrl),
	.cout());
defparam \sink_ready_ctrl~2 .lut_mask = 16'hFEFF;
defparam \sink_ready_ctrl~2 .sum_lutc_input = "datac";

dffeas stall_reg(
	.clk(clk),
	.d(\stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stall_reg1),
	.prn(vcc));
defparam stall_reg.is_wysiwyg = "true";
defparam stall_reg.power_up = "low";

cycloneive_lcell_comb \sink_ready_ctrl~0 (
	.dataa(\ready_FIFO|fifo_array[5][0]~q ),
	.datab(\ready_FIFO|fifo_array[4][0]~q ),
	.datac(gnd),
	.datad(\ready_FIFO|rd_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\sink_ready_ctrl~0_combout ),
	.cout());
defparam \sink_ready_ctrl~0 .lut_mask = 16'hAACC;
defparam \sink_ready_ctrl~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready_ctrl~1 (
	.dataa(\sink_ready_ctrl~0_combout ),
	.datab(\ready_FIFO|rd_addr_ptr[2]~q ),
	.datac(gnd),
	.datad(\ready_FIFO|rd_addr_ptr[1]~q ),
	.cin(gnd),
	.combout(\sink_ready_ctrl~1_combout ),
	.cout());
defparam \sink_ready_ctrl~1 .lut_mask = 16'hEEFF;
defparam \sink_ready_ctrl~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \stall_reg~0 (
	.dataa(dffe_af),
	.datab(gnd),
	.datac(dffe_nae),
	.datad(reset_n),
	.cin(gnd),
	.combout(\stall_reg~0_combout ),
	.cout());
defparam \stall_reg~0 .lut_mask = 16'hAFFF;
defparam \stall_reg~0 .sum_lutc_input = "datac";

endmodule

module CIC_auk_dspip_avalon_streaming_small_fifo (
	dffe_nae,
	fifo_array_0_5,
	fifo_array_0_4,
	rd_addr_ptr_2,
	dffe_af,
	rd_addr_ptr_0,
	rd_addr_ptr_1,
	Equal2,
	Mux0,
	stall_reg,
	usedw_process,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	dffe_nae;
output 	fifo_array_0_5;
output 	fifo_array_0_4;
output 	rd_addr_ptr_2;
input 	dffe_af;
output 	rd_addr_ptr_0;
output 	rd_addr_ptr_1;
output 	Equal2;
output 	Mux0;
input 	stall_reg;
output 	usedw_process;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_addr_ptr~2_combout ;
wire \fifo_usedw[2]~0_combout ;
wire \fifo_usedw[0]~2_combout ;
wire \fifo_usedw[0]~3_combout ;
wire \fifo_usedw[0]~q ;
wire \usedw_process~2_combout ;
wire \Add2~1_combout ;
wire \fifo_usedw[1]~4_combout ;
wire \fifo_usedw[1]~q ;
wire \Add2~0_combout ;
wire \fifo_usedw[2]~1_combout ;
wire \fifo_usedw[2]~q ;
wire \usedw_process~1_combout ;
wire \wr_addr_ptr[0]~1_combout ;
wire \wr_addr_ptr[0]~q ;
wire \wr_addr_ptr~3_combout ;
wire \wr_addr_ptr[2]~q ;
wire \wr_addr_ptr~0_combout ;
wire \wr_addr_ptr[1]~q ;
wire \Decoder0~0_combout ;
wire \fifo_array~0_combout ;
wire \fifo_array~1_combout ;
wire \rd_addr_ptr~3_combout ;
wire \rd_addr_ptr[1]~5_combout ;
wire \rd_addr_ptr~2_combout ;
wire \rd_addr_ptr~4_combout ;
wire \Decoder0~1_combout ;
wire \Decoder0~2_combout ;
wire \fifo_array~2_combout ;
wire \fifo_array[2][0]~q ;
wire \fifo_array~3_combout ;
wire \fifo_array[1][0]~q ;
wire \fifo_array~4_combout ;
wire \fifo_array[0][0]~q ;
wire \Mux0~0_combout ;
wire \fifo_array~5_combout ;
wire \fifo_array[3][0]~q ;


dffeas \fifo_array[5][0] (
	.clk(clock),
	.d(\fifo_array~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_array_0_5),
	.prn(vcc));
defparam \fifo_array[5][0] .is_wysiwyg = "true";
defparam \fifo_array[5][0] .power_up = "low";

dffeas \fifo_array[4][0] (
	.clk(clock),
	.d(\fifo_array~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_array_0_4),
	.prn(vcc));
defparam \fifo_array[4][0] .is_wysiwyg = "true";
defparam \fifo_array[4][0] .power_up = "low";

dffeas \rd_addr_ptr[2] (
	.clk(clock),
	.d(\rd_addr_ptr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\rd_addr_ptr[1]~5_combout ),
	.q(rd_addr_ptr_2),
	.prn(vcc));
defparam \rd_addr_ptr[2] .is_wysiwyg = "true";
defparam \rd_addr_ptr[2] .power_up = "low";

dffeas \rd_addr_ptr[0] (
	.clk(clock),
	.d(\rd_addr_ptr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_addr_ptr[1]~5_combout ),
	.q(rd_addr_ptr_0),
	.prn(vcc));
defparam \rd_addr_ptr[0] .is_wysiwyg = "true";
defparam \rd_addr_ptr[0] .power_up = "low";

dffeas \rd_addr_ptr[1] (
	.clk(clock),
	.d(\rd_addr_ptr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_addr_ptr[1]~5_combout ),
	.q(rd_addr_ptr_1),
	.prn(vcc));
defparam \rd_addr_ptr[1] .is_wysiwyg = "true";
defparam \rd_addr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(gnd),
	.datab(\fifo_usedw[2]~q ),
	.datac(\fifo_usedw[0]~q ),
	.datad(\fifo_usedw[1]~q ),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h3FFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\fifo_array[2][0]~q ),
	.datab(rd_addr_ptr_1),
	.datac(\Mux0~0_combout ),
	.datad(\fifo_array[3][0]~q ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_process~0 (
	.dataa(dffe_nae),
	.datab(gnd),
	.datac(gnd),
	.datad(dffe_af),
	.cin(gnd),
	.combout(usedw_process),
	.cout());
defparam \usedw_process~0 .lut_mask = 16'hAAFF;
defparam \usedw_process~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_addr_ptr~2 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\wr_addr_ptr~2_combout ),
	.cout());
defparam \wr_addr_ptr~2 .lut_mask = 16'hAAFF;
defparam \wr_addr_ptr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_usedw[2]~0 (
	.dataa(usedw_process),
	.datab(\usedw_process~1_combout ),
	.datac(Equal2),
	.datad(reset_n),
	.cin(gnd),
	.combout(\fifo_usedw[2]~0_combout ),
	.cout());
defparam \fifo_usedw[2]~0 .lut_mask = 16'h6FFF;
defparam \fifo_usedw[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_usedw[0]~2 (
	.dataa(\fifo_usedw[0]~q ),
	.datab(Equal2),
	.datac(usedw_process),
	.datad(\usedw_process~1_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[0]~2_combout ),
	.cout());
defparam \fifo_usedw[0]~2 .lut_mask = 16'h6996;
defparam \fifo_usedw[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_usedw[0]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(reset_n),
	.datad(\fifo_usedw[0]~2_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[0]~3_combout ),
	.cout());
defparam \fifo_usedw[0]~3 .lut_mask = 16'hFFF0;
defparam \fifo_usedw[0]~3 .sum_lutc_input = "datac";

dffeas \fifo_usedw[0] (
	.clk(clock),
	.d(\fifo_usedw[0]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[0]~q ),
	.prn(vcc));
defparam \fifo_usedw[0] .is_wysiwyg = "true";
defparam \fifo_usedw[0] .power_up = "low";

cycloneive_lcell_comb \usedw_process~2 (
	.dataa(dffe_af),
	.datab(gnd),
	.datac(dffe_nae),
	.datad(\usedw_process~1_combout ),
	.cin(gnd),
	.combout(\usedw_process~2_combout ),
	.cout());
defparam \usedw_process~2 .lut_mask = 16'hAFFF;
defparam \usedw_process~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add2~1 (
	.dataa(\fifo_usedw[0]~q ),
	.datab(\fifo_usedw[1]~q ),
	.datac(\usedw_process~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h9696;
defparam \Add2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_usedw[1]~4 (
	.dataa(\fifo_usedw[1]~q ),
	.datab(reset_n),
	.datac(\fifo_usedw[2]~0_combout ),
	.datad(\Add2~1_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[1]~4_combout ),
	.cout());
defparam \fifo_usedw[1]~4 .lut_mask = 16'hACFF;
defparam \fifo_usedw[1]~4 .sum_lutc_input = "datac";

dffeas \fifo_usedw[1] (
	.clk(clock),
	.d(\fifo_usedw[1]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[1]~q ),
	.prn(vcc));
defparam \fifo_usedw[1] .is_wysiwyg = "true";
defparam \fifo_usedw[1] .power_up = "low";

cycloneive_lcell_comb \Add2~0 (
	.dataa(\fifo_usedw[0]~q ),
	.datab(\fifo_usedw[1]~q ),
	.datac(\usedw_process~2_combout ),
	.datad(\fifo_usedw[2]~q ),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h6996;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_usedw[2]~1 (
	.dataa(\fifo_usedw[2]~q ),
	.datab(reset_n),
	.datac(\fifo_usedw[2]~0_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[2]~1_combout ),
	.cout());
defparam \fifo_usedw[2]~1 .lut_mask = 16'hACFF;
defparam \fifo_usedw[2]~1 .sum_lutc_input = "datac";

dffeas \fifo_usedw[2] (
	.clk(clock),
	.d(\fifo_usedw[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[2]~q ),
	.prn(vcc));
defparam \fifo_usedw[2] .is_wysiwyg = "true";
defparam \fifo_usedw[2] .power_up = "low";

cycloneive_lcell_comb \usedw_process~1 (
	.dataa(stall_reg),
	.datab(\fifo_usedw[2]~q ),
	.datac(\fifo_usedw[1]~q ),
	.datad(\fifo_usedw[0]~q ),
	.cin(gnd),
	.combout(\usedw_process~1_combout ),
	.cout());
defparam \usedw_process~1 .lut_mask = 16'hFEFF;
defparam \usedw_process~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_addr_ptr[0]~1 (
	.dataa(reset_n),
	.datab(\usedw_process~1_combout ),
	.datac(usedw_process),
	.datad(Equal2),
	.cin(gnd),
	.combout(\wr_addr_ptr[0]~1_combout ),
	.cout());
defparam \wr_addr_ptr[0]~1 .lut_mask = 16'h7FFF;
defparam \wr_addr_ptr[0]~1 .sum_lutc_input = "datac";

dffeas \wr_addr_ptr[0] (
	.clk(clock),
	.d(\wr_addr_ptr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_ptr[0]~1_combout ),
	.q(\wr_addr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[0] .is_wysiwyg = "true";
defparam \wr_addr_ptr[0] .power_up = "low";

cycloneive_lcell_comb \wr_addr_ptr~3 (
	.dataa(\wr_addr_ptr[1]~q ),
	.datab(gnd),
	.datac(\wr_addr_ptr[2]~q ),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\wr_addr_ptr~3_combout ),
	.cout());
defparam \wr_addr_ptr~3 .lut_mask = 16'hAFFA;
defparam \wr_addr_ptr~3 .sum_lutc_input = "datac";

dffeas \wr_addr_ptr[2] (
	.clk(clock),
	.d(\wr_addr_ptr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\wr_addr_ptr[0]~1_combout ),
	.q(\wr_addr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[2] .is_wysiwyg = "true";
defparam \wr_addr_ptr[2] .power_up = "low";

cycloneive_lcell_comb \wr_addr_ptr~0 (
	.dataa(reset_n),
	.datab(\wr_addr_ptr[1]~q ),
	.datac(\wr_addr_ptr[2]~q ),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\wr_addr_ptr~0_combout ),
	.cout());
defparam \wr_addr_ptr~0 .lut_mask = 16'hBFEF;
defparam \wr_addr_ptr~0 .sum_lutc_input = "datac";

dffeas \wr_addr_ptr[1] (
	.clk(clock),
	.d(\wr_addr_ptr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_ptr[0]~1_combout ),
	.q(\wr_addr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[1] .is_wysiwyg = "true";
defparam \wr_addr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \Decoder0~0 (
	.dataa(usedw_process),
	.datab(Equal2),
	.datac(\wr_addr_ptr[1]~q ),
	.datad(\usedw_process~1_combout ),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
defparam \Decoder0~0 .lut_mask = 16'h7FFF;
defparam \Decoder0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_array~0 (
	.dataa(fifo_array_0_5),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[0]~q ),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\fifo_array~0_combout ),
	.cout());
defparam \fifo_array~0 .lut_mask = 16'hFFFE;
defparam \fifo_array~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_array~1 (
	.dataa(fifo_array_0_4),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[2]~q ),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\fifo_array~1_combout ),
	.cout());
defparam \fifo_array~1 .lut_mask = 16'hFEFF;
defparam \fifo_array~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_ptr~3 (
	.dataa(rd_addr_ptr_1),
	.datab(gnd),
	.datac(rd_addr_ptr_2),
	.datad(rd_addr_ptr_0),
	.cin(gnd),
	.combout(\rd_addr_ptr~3_combout ),
	.cout());
defparam \rd_addr_ptr~3 .lut_mask = 16'hAFFA;
defparam \rd_addr_ptr~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_ptr[1]~5 (
	.dataa(dffe_nae),
	.datab(dffe_af),
	.datac(reset_n),
	.datad(Equal2),
	.cin(gnd),
	.combout(\rd_addr_ptr[1]~5_combout ),
	.cout());
defparam \rd_addr_ptr[1]~5 .lut_mask = 16'hBFFF;
defparam \rd_addr_ptr[1]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_ptr~2 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(rd_addr_ptr_0),
	.cin(gnd),
	.combout(\rd_addr_ptr~2_combout ),
	.cout());
defparam \rd_addr_ptr~2 .lut_mask = 16'hAAFF;
defparam \rd_addr_ptr~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_addr_ptr~4 (
	.dataa(reset_n),
	.datab(rd_addr_ptr_1),
	.datac(rd_addr_ptr_2),
	.datad(rd_addr_ptr_0),
	.cin(gnd),
	.combout(\rd_addr_ptr~4_combout ),
	.cout());
defparam \rd_addr_ptr~4 .lut_mask = 16'hBFEF;
defparam \rd_addr_ptr~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~1 (
	.dataa(\wr_addr_ptr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
defparam \Decoder0~1 .lut_mask = 16'hAAFF;
defparam \Decoder0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Decoder0~2 (
	.dataa(\Decoder0~1_combout ),
	.datab(usedw_process),
	.datac(Equal2),
	.datad(\usedw_process~1_combout ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
defparam \Decoder0~2 .lut_mask = 16'hBFFF;
defparam \Decoder0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_array~2 (
	.dataa(\fifo_array[2][0]~q ),
	.datab(\Decoder0~2_combout ),
	.datac(gnd),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\fifo_array~2_combout ),
	.cout());
defparam \fifo_array~2 .lut_mask = 16'hEEFF;
defparam \fifo_array~2 .sum_lutc_input = "datac";

dffeas \fifo_array[2][0] (
	.clk(clock),
	.d(\fifo_array~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[2][0]~q ),
	.prn(vcc));
defparam \fifo_array[2][0] .is_wysiwyg = "true";
defparam \fifo_array[2][0] .power_up = "low";

cycloneive_lcell_comb \fifo_array~3 (
	.dataa(\fifo_array[1][0]~q ),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[0]~q ),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\fifo_array~3_combout ),
	.cout());
defparam \fifo_array~3 .lut_mask = 16'hFEFF;
defparam \fifo_array~3 .sum_lutc_input = "datac";

dffeas \fifo_array[1][0] (
	.clk(clock),
	.d(\fifo_array~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[1][0]~q ),
	.prn(vcc));
defparam \fifo_array[1][0] .is_wysiwyg = "true";
defparam \fifo_array[1][0] .power_up = "low";

cycloneive_lcell_comb \fifo_array~4 (
	.dataa(\fifo_array[0][0]~q ),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[0]~q ),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\fifo_array~4_combout ),
	.cout());
defparam \fifo_array~4 .lut_mask = 16'hEFFF;
defparam \fifo_array~4 .sum_lutc_input = "datac";

dffeas \fifo_array[0][0] (
	.clk(clock),
	.d(\fifo_array~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[0][0]~q ),
	.prn(vcc));
defparam \fifo_array[0][0] .is_wysiwyg = "true";
defparam \fifo_array[0][0] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(rd_addr_ptr_1),
	.datab(\fifo_array[1][0]~q ),
	.datac(rd_addr_ptr_0),
	.datad(\fifo_array[0][0]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_array~5 (
	.dataa(\fifo_array[3][0]~q ),
	.datab(\wr_addr_ptr[0]~q ),
	.datac(\Decoder0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_array~5_combout ),
	.cout());
defparam \fifo_array~5 .lut_mask = 16'hFEFE;
defparam \fifo_array~5 .sum_lutc_input = "datac";

dffeas \fifo_array[3][0] (
	.clk(clock),
	.d(\fifo_array~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[3][0]~q ),
	.prn(vcc));
defparam \fifo_array[3][0] .is_wysiwyg = "true";
defparam \fifo_array[3][0] .power_up = "low";

endmodule

module CIC_auk_dspip_avalon_streaming_sink (
	full_dff,
	dffe_nae,
	dffe_af,
	data,
	sink_ready_ctrl,
	usedw_process,
	GND_port,
	clk,
	in_valid,
	reset_n,
	at_sink_data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	dffe_nae;
input 	dffe_af;
output 	[255:0] data;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	GND_port;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	[255:0] at_sink_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_17 sink_FIFO(
	.full_dff(full_dff),
	.dffe_nae(dffe_nae),
	.dffe_af(dffe_af),
	.q({q_unconnected_wire_257,q_unconnected_wire_256,data[255],data[254],data[253],data[252],data[251],data[250],data[249],data[248],data[247],data[246],data[245],data[244],q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,data[239],data[238],data[237],data[236],data[235],data[234],data[233],data[232],data[231],data[230],data[229],data[228],q_unconnected_wire_227,
q_unconnected_wire_226,q_unconnected_wire_225,q_unconnected_wire_224,data[223],data[222],data[221],data[220],data[219],data[218],data[217],data[216],data[215],data[214],data[213],data[212],q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,data[207],data[206],data[205],data[204],data[203],data[202],data[201],data[200],data[199],data[198],data[197],data[196],
q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,data[191],data[190],data[189],data[188],data[187],data[186],data[185],data[184],data[183],data[182],data[181],data[180],q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,data[175],data[174],data[173],data[172],data[171],data[170],data[169],data[168],
data[167],data[166],data[165],data[164],q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,data[159],data[158],data[157],data[156],data[155],data[154],data[153],data[152],data[151],data[150],data[149],data[148],q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,data[143],data[142],data[141],data[140],
data[139],data[138],data[137],data[136],data[135],data[134],data[133],data[132],q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,data[127],data[126],data[125],data[124],data[123],data[122],data[121],data[120],data[119],data[118],data[117],data[116],q_unconnected_wire_115,q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,
data[111],data[110],data[109],data[108],data[107],data[106],data[105],data[104],data[103],data[102],data[101],data[100],q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,data[95],data[94],data[93],data[92],data[91],data[90],data[89],data[88],data[87],data[86],data[85],data[84],q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,
q_unconnected_wire_80,data[79],data[78],data[77],data[76],data[75],data[74],data[73],data[72],data[71],data[70],data[69],data[68],q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,data[63],data[62],data[61],data[60],data[59],data[58],data[57],data[56],data[55],data[54],data[53],data[52],q_unconnected_wire_51,q_unconnected_wire_50,
q_unconnected_wire_49,q_unconnected_wire_48,data[47],data[46],data[45],data[44],data[43],data[42],data[41],data[40],data[39],data[38],data[37],data[36],q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],q_unconnected_wire_19,
q_unconnected_wire_18,q_unconnected_wire_17,q_unconnected_wire_16,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.sink_ready_ctrl(sink_ready_ctrl),
	.usedw_process(usedw_process),
	.GND_port(GND_port),
	.clock(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.data({gnd,gnd,at_sink_data[255],at_sink_data[254],at_sink_data[253],at_sink_data[252],at_sink_data[251],at_sink_data[250],at_sink_data[249],at_sink_data[248],at_sink_data[247],at_sink_data[246],at_sink_data[245],at_sink_data[244],gnd,gnd,gnd,gnd,at_sink_data[239],at_sink_data[238],at_sink_data[237],at_sink_data[236],at_sink_data[235],at_sink_data[234],at_sink_data[233],
at_sink_data[232],at_sink_data[231],at_sink_data[230],at_sink_data[229],at_sink_data[228],gnd,gnd,gnd,gnd,at_sink_data[223],at_sink_data[222],at_sink_data[221],at_sink_data[220],at_sink_data[219],at_sink_data[218],at_sink_data[217],at_sink_data[216],at_sink_data[215],at_sink_data[214],at_sink_data[213],at_sink_data[212],gnd,gnd,gnd,gnd,at_sink_data[207],at_sink_data[206],
at_sink_data[205],at_sink_data[204],at_sink_data[203],at_sink_data[202],at_sink_data[201],at_sink_data[200],at_sink_data[199],at_sink_data[198],at_sink_data[197],at_sink_data[196],gnd,gnd,gnd,gnd,at_sink_data[191],at_sink_data[190],at_sink_data[189],at_sink_data[188],at_sink_data[187],at_sink_data[186],at_sink_data[185],at_sink_data[184],at_sink_data[183],at_sink_data[182],
at_sink_data[181],at_sink_data[180],gnd,gnd,gnd,gnd,at_sink_data[175],at_sink_data[174],at_sink_data[173],at_sink_data[172],at_sink_data[171],at_sink_data[170],at_sink_data[169],at_sink_data[168],at_sink_data[167],at_sink_data[166],at_sink_data[165],at_sink_data[164],gnd,gnd,gnd,gnd,at_sink_data[159],at_sink_data[158],at_sink_data[157],at_sink_data[156],at_sink_data[155],
at_sink_data[154],at_sink_data[153],at_sink_data[152],at_sink_data[151],at_sink_data[150],at_sink_data[149],at_sink_data[148],gnd,gnd,gnd,gnd,at_sink_data[143],at_sink_data[142],at_sink_data[141],at_sink_data[140],at_sink_data[139],at_sink_data[138],at_sink_data[137],at_sink_data[136],at_sink_data[135],at_sink_data[134],at_sink_data[133],at_sink_data[132],gnd,gnd,gnd,gnd,
at_sink_data[127],at_sink_data[126],at_sink_data[125],at_sink_data[124],at_sink_data[123],at_sink_data[122],at_sink_data[121],at_sink_data[120],at_sink_data[119],at_sink_data[118],at_sink_data[117],at_sink_data[116],gnd,gnd,gnd,gnd,at_sink_data[111],at_sink_data[110],at_sink_data[109],at_sink_data[108],at_sink_data[107],at_sink_data[106],at_sink_data[105],at_sink_data[104],
at_sink_data[103],at_sink_data[102],at_sink_data[101],at_sink_data[100],gnd,gnd,gnd,gnd,at_sink_data[95],at_sink_data[94],at_sink_data[93],at_sink_data[92],at_sink_data[91],at_sink_data[90],at_sink_data[89],at_sink_data[88],at_sink_data[87],at_sink_data[86],at_sink_data[85],at_sink_data[84],gnd,gnd,gnd,gnd,at_sink_data[79],at_sink_data[78],at_sink_data[77],
at_sink_data[76],at_sink_data[75],at_sink_data[74],at_sink_data[73],at_sink_data[72],at_sink_data[71],at_sink_data[70],at_sink_data[69],at_sink_data[68],gnd,gnd,gnd,gnd,at_sink_data[63],at_sink_data[62],at_sink_data[61],at_sink_data[60],at_sink_data[59],at_sink_data[58],at_sink_data[57],at_sink_data[56],at_sink_data[55],at_sink_data[54],at_sink_data[53],
at_sink_data[52],gnd,gnd,gnd,gnd,at_sink_data[47],at_sink_data[46],at_sink_data[45],at_sink_data[44],at_sink_data[43],at_sink_data[42],at_sink_data[41],at_sink_data[40],at_sink_data[39],at_sink_data[38],at_sink_data[37],at_sink_data[36],gnd,gnd,gnd,gnd,at_sink_data[31],at_sink_data[30],at_sink_data[29],at_sink_data[28],at_sink_data[27],at_sink_data[26],
at_sink_data[25],at_sink_data[24],at_sink_data[23],at_sink_data[22],at_sink_data[21],at_sink_data[20],gnd,gnd,gnd,gnd,at_sink_data[15],at_sink_data[14],at_sink_data[13],at_sink_data[12],at_sink_data[11],at_sink_data[10],at_sink_data[9],at_sink_data[8],at_sink_data[7],at_sink_data[6],at_sink_data[5],at_sink_data[4],gnd,gnd,gnd,gnd}));

endmodule

module CIC_scfifo_17 (
	full_dff,
	dffe_nae,
	dffe_af,
	q,
	sink_ready_ctrl,
	usedw_process,
	GND_port,
	clock,
	in_valid,
	reset_n,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	dffe_nae;
input 	dffe_af;
output 	[257:0] q;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;
input 	[257:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_6h71 auto_generated(
	.full_dff(full_dff),
	.dffe_nae1(dffe_nae),
	.dffe_af(dffe_af),
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q[255],q[254],q[253],q[252],q[251],q[250],q[249],q[248],q[247],q[246],q[245],q[244],q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q[239],q[238],q[237],q[236],q[235],q[234],q[233],q[232],q[231],q[230],q[229],q[228],q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,q_unconnected_wire_224,q[223],q[222],q[221],q[220],q[219],q[218],q[217],q[216],q[215],q[214],q[213],q[212],
q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q[207],q[206],q[205],q[204],q[203],q[202],q[201],q[200],q[199],q[198],q[197],q[196],q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,q[191],q[190],q[189],q[188],q[187],q[186],q[185],q[184],q[183],q[182],q[181],q[180],q_unconnected_wire_179,q_unconnected_wire_178,
q_unconnected_wire_177,q_unconnected_wire_176,q[175],q[174],q[173],q[172],q[171],q[170],q[169],q[168],q[167],q[166],q[165],q[164],q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q[159],q[158],q[157],q[156],q[155],q[154],q[153],q[152],q[151],q[150],q[149],q[148],q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q[143],q[142],q[141],q[140],q[139],q[138],q[137],q[136],q[135],q[134],q[133],q[132],
q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q[127],q[126],q[125],q[124],q[123],q[122],q[121],q[120],q[119],q[118],q[117],q[116],q_unconnected_wire_115,q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q[111],q[110],q[109],q[108],q[107],q[106],q[105],q[104],q[103],q[102],q[101],q[100],q_unconnected_wire_99,q_unconnected_wire_98,
q_unconnected_wire_97,q_unconnected_wire_96,q[95],q[94],q[93],q[92],q[91],q[90],q[89],q[88],q[87],q[86],q[85],q[84],q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,q[79],q[78],q[77],q[76],q[75],q[74],q[73],q[72],q[71],q[70],q[69],q[68],q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q[63],q[62],q[61],q[60],q[59],q[58],q[57],q[56],q[55],q[54],q[53],q[52],
q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q[47],q[46],q[45],q[44],q[43],q[42],q[41],q[40],q[39],q[38],q[37],q[36],q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q_unconnected_wire_19,q_unconnected_wire_18,q_unconnected_wire_17,
q_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.sink_ready_ctrl(sink_ready_ctrl),
	.usedw_process(usedw_process),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.data({gnd,gnd,data[255],data[254],data[253],data[252],data[251],data[250],data[249],data[248],data[247],data[246],data[245],data[244],gnd,gnd,gnd,gnd,data[239],data[238],data[237],data[236],data[235],data[234],data[233],data[232],data[231],data[230],data[229],data[228],gnd,gnd,gnd,gnd,data[223],data[222],data[221],data[220],data[219],data[218],data[217],data[216],data[215],data[214],data[213],data[212],gnd,gnd,gnd,gnd,data[207],data[206],data[205],data[204],data[203],data[202],data[201],data[200],data[199],data[198],data[197],data[196],gnd,gnd,gnd,gnd,data[191],data[190],
data[189],data[188],data[187],data[186],data[185],data[184],data[183],data[182],data[181],data[180],gnd,gnd,gnd,gnd,data[175],data[174],data[173],data[172],data[171],data[170],data[169],data[168],data[167],data[166],data[165],data[164],gnd,gnd,gnd,gnd,data[159],data[158],data[157],data[156],data[155],data[154],data[153],data[152],data[151],data[150],data[149],data[148],gnd,gnd,gnd,gnd,data[143],data[142],data[141],data[140],data[139],data[138],data[137],data[136],data[135],data[134],data[133],data[132],gnd,gnd,gnd,gnd,data[127],data[126],data[125],data[124],data[123],data[122],
data[121],data[120],data[119],data[118],data[117],data[116],gnd,gnd,gnd,gnd,data[111],data[110],data[109],data[108],data[107],data[106],data[105],data[104],data[103],data[102],data[101],data[100],gnd,gnd,gnd,gnd,data[95],data[94],data[93],data[92],data[91],data[90],data[89],data[88],data[87],data[86],data[85],data[84],gnd,gnd,gnd,gnd,data[79],data[78],data[77],data[76],data[75],data[74],data[73],data[72],data[71],data[70],data[69],data[68],gnd,gnd,gnd,gnd,data[63],data[62],data[61],data[60],data[59],data[58],data[57],data[56],data[55],data[54],
data[53],data[52],gnd,gnd,gnd,gnd,data[47],data[46],data[45],data[44],data[43],data[42],data[41],data[40],data[39],data[38],data[37],data[36],gnd,gnd,gnd,gnd,data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],gnd,gnd,gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],gnd,gnd,gnd,gnd}));

endmodule

module CIC_scfifo_6h71 (
	full_dff,
	dffe_nae1,
	dffe_af,
	q,
	sink_ready_ctrl,
	usedw_process,
	GND_port,
	clock,
	in_valid,
	reset_n,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	dffe_nae1;
input 	dffe_af;
output 	[257:0] q;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;
input 	[257:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \dffe_nae~2_combout ;
wire \dffe_nae~3_combout ;
wire \dffe_nae~4_combout ;


CIC_a_dpfifo_nmv dpfifo(
	.full_dff1(full_dff),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.dffe_nae(dffe_nae1),
	.dffe_af(dffe_af),
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q[255],q[254],q[253],q[252],q[251],q[250],q[249],q[248],q[247],q[246],q[245],q[244],q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q[239],q[238],q[237],q[236],q[235],q[234],q[233],q[232],q[231],q[230],q[229],q[228],q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,q_unconnected_wire_224,q[223],q[222],q[221],q[220],q[219],q[218],q[217],q[216],q[215],q[214],q[213],q[212],
q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q[207],q[206],q[205],q[204],q[203],q[202],q[201],q[200],q[199],q[198],q[197],q[196],q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,q[191],q[190],q[189],q[188],q[187],q[186],q[185],q[184],q[183],q[182],q[181],q[180],q_unconnected_wire_179,q_unconnected_wire_178,
q_unconnected_wire_177,q_unconnected_wire_176,q[175],q[174],q[173],q[172],q[171],q[170],q[169],q[168],q[167],q[166],q[165],q[164],q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q[159],q[158],q[157],q[156],q[155],q[154],q[153],q[152],q[151],q[150],q[149],q[148],q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q[143],q[142],q[141],q[140],q[139],q[138],q[137],q[136],q[135],q[134],q[133],q[132],
q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q[127],q[126],q[125],q[124],q[123],q[122],q[121],q[120],q[119],q[118],q[117],q[116],q_unconnected_wire_115,q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q[111],q[110],q[109],q[108],q[107],q[106],q[105],q[104],q[103],q[102],q[101],q[100],q_unconnected_wire_99,q_unconnected_wire_98,
q_unconnected_wire_97,q_unconnected_wire_96,q[95],q[94],q[93],q[92],q[91],q[90],q[89],q[88],q[87],q[86],q[85],q[84],q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,q[79],q[78],q[77],q[76],q[75],q[74],q[73],q[72],q[71],q[70],q[69],q[68],q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q[63],q[62],q[61],q[60],q[59],q[58],q[57],q[56],q[55],q[54],q[53],q[52],
q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q[47],q[46],q[45],q[44],q[43],q[42],q[41],q[40],q[39],q[38],q[37],q[36],q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q_unconnected_wire_19,q_unconnected_wire_18,q_unconnected_wire_17,
q_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q_unconnected_wire_3,q_unconnected_wire_2,q_unconnected_wire_1,q_unconnected_wire_0}),
	.sink_ready_ctrl(sink_ready_ctrl),
	.usedw_process(usedw_process),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.data({gnd,gnd,data[255],data[254],data[253],data[252],data[251],data[250],data[249],data[248],data[247],data[246],data[245],data[244],gnd,gnd,gnd,gnd,data[239],data[238],data[237],data[236],data[235],data[234],data[233],data[232],data[231],data[230],data[229],data[228],gnd,gnd,gnd,gnd,data[223],data[222],data[221],data[220],data[219],data[218],data[217],data[216],data[215],data[214],data[213],data[212],gnd,gnd,gnd,gnd,data[207],data[206],data[205],data[204],data[203],data[202],data[201],data[200],data[199],data[198],data[197],data[196],gnd,gnd,gnd,gnd,data[191],data[190],
data[189],data[188],data[187],data[186],data[185],data[184],data[183],data[182],data[181],data[180],gnd,gnd,gnd,gnd,data[175],data[174],data[173],data[172],data[171],data[170],data[169],data[168],data[167],data[166],data[165],data[164],gnd,gnd,gnd,gnd,data[159],data[158],data[157],data[156],data[155],data[154],data[153],data[152],data[151],data[150],data[149],data[148],gnd,gnd,gnd,gnd,data[143],data[142],data[141],data[140],data[139],data[138],data[137],data[136],data[135],data[134],data[133],data[132],gnd,gnd,gnd,gnd,data[127],data[126],data[125],data[124],data[123],data[122],
data[121],data[120],data[119],data[118],data[117],data[116],gnd,gnd,gnd,gnd,data[111],data[110],data[109],data[108],data[107],data[106],data[105],data[104],data[103],data[102],data[101],data[100],gnd,gnd,gnd,gnd,data[95],data[94],data[93],data[92],data[91],data[90],data[89],data[88],data[87],data[86],data[85],data[84],gnd,gnd,gnd,gnd,data[79],data[78],data[77],data[76],data[75],data[74],data[73],data[72],data[71],data[70],data[69],data[68],gnd,gnd,gnd,gnd,data[63],data[62],data[61],data[60],data[59],data[58],data[57],data[56],data[55],data[54],
data[53],data[52],gnd,gnd,gnd,gnd,data[47],data[46],data[45],data[44],data[43],data[42],data[41],data[40],data[39],data[38],data[37],data[36],gnd,gnd,gnd,gnd,data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],gnd,gnd,gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],gnd,gnd,gnd,gnd}));

dffeas dffe_nae(
	.clk(clock),
	.d(\dffe_nae~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_nae1),
	.prn(vcc));
defparam dffe_nae.is_wysiwyg = "true";
defparam dffe_nae.power_up = "low";

cycloneive_lcell_comb \dffe_nae~2 (
	.dataa(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(dffe_nae1),
	.datad(gnd),
	.cin(gnd),
	.combout(\dffe_nae~2_combout ),
	.cout());
defparam \dffe_nae~2 .lut_mask = 16'hFEFE;
defparam \dffe_nae~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe_nae~3 (
	.dataa(in_valid),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datac(dffe_nae1),
	.datad(\dffe_nae~2_combout ),
	.cin(gnd),
	.combout(\dffe_nae~3_combout ),
	.cout());
defparam \dffe_nae~3 .lut_mask = 16'h6996;
defparam \dffe_nae~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe_nae~4 (
	.dataa(dffe_nae1),
	.datab(dffe_af),
	.datac(sink_ready_ctrl),
	.datad(\dffe_nae~3_combout ),
	.cin(gnd),
	.combout(\dffe_nae~4_combout ),
	.cout());
defparam \dffe_nae~4 .lut_mask = 16'hDFEF;
defparam \dffe_nae~4 .sum_lutc_input = "datac";

endmodule

module CIC_a_dpfifo_nmv (
	full_dff1,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	dffe_nae,
	dffe_af,
	q,
	sink_ready_ctrl,
	usedw_process,
	GND_port,
	clock,
	in_valid,
	reset_n,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	dffe_nae;
input 	dffe_af;
output 	[257:0] q;
input 	sink_ready_ctrl;
input 	usedw_process;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;
input 	[257:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \_~0_combout ;
wire \empty_dff~2_combout ;
wire \usedw_is_0_dff~q ;
wire \valid_wreq~combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \empty_dff~1_combout ;
wire \empty_dff~q ;
wire \valid_rreq~combout ;
wire \_~1_combout ;


CIC_cntr_s9b wr_ptr(
	.full_dff(full_dff1),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n));

CIC_cntr_8a7 usedw_counter(
	.full_dff(full_dff1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.valid_rreq(\valid_rreq~combout ),
	.updown(\valid_wreq~combout ),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n));

CIC_cntr_r9b rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.valid_rreq(\valid_rreq~combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_1bh1 FIFOram(
	.q_b({q_b_unconnected_wire_257,q_b_unconnected_wire_256,q[255],q[254],q[253],q[252],q[251],q[250],q[249],q[248],q[247],q[246],q[245],q[244],q_b_unconnected_wire_243,q_b_unconnected_wire_242,q_b_unconnected_wire_241,q_b_unconnected_wire_240,q[239],q[238],q[237],q[236],q[235],q[234],q[233],q[232],q[231],q[230],q[229],q[228],q_b_unconnected_wire_227,q_b_unconnected_wire_226,q_b_unconnected_wire_225,
q_b_unconnected_wire_224,q[223],q[222],q[221],q[220],q[219],q[218],q[217],q[216],q[215],q[214],q[213],q[212],q_b_unconnected_wire_211,q_b_unconnected_wire_210,q_b_unconnected_wire_209,q_b_unconnected_wire_208,q[207],q[206],q[205],q[204],q[203],q[202],q[201],q[200],q[199],q[198],q[197],q[196],q_b_unconnected_wire_195,q_b_unconnected_wire_194,q_b_unconnected_wire_193,q_b_unconnected_wire_192,q[191],q[190],q[189],q[188],q[187],q[186],q[185],q[184],q[183],q[182],q[181],q[180],
q_b_unconnected_wire_179,q_b_unconnected_wire_178,q_b_unconnected_wire_177,q_b_unconnected_wire_176,q[175],q[174],q[173],q[172],q[171],q[170],q[169],q[168],q[167],q[166],q[165],q[164],q_b_unconnected_wire_163,q_b_unconnected_wire_162,q_b_unconnected_wire_161,q_b_unconnected_wire_160,q[159],q[158],q[157],q[156],q[155],q[154],q[153],q[152],q[151],q[150],q[149],q[148],q_b_unconnected_wire_147,
q_b_unconnected_wire_146,q_b_unconnected_wire_145,q_b_unconnected_wire_144,q[143],q[142],q[141],q[140],q[139],q[138],q[137],q[136],q[135],q[134],q[133],q[132],q_b_unconnected_wire_131,q_b_unconnected_wire_130,q_b_unconnected_wire_129,q_b_unconnected_wire_128,q[127],q[126],q[125],q[124],q[123],q[122],q[121],q[120],q[119],q[118],q[117],q[116],q_b_unconnected_wire_115,q_b_unconnected_wire_114,
q_b_unconnected_wire_113,q_b_unconnected_wire_112,q[111],q[110],q[109],q[108],q[107],q[106],q[105],q[104],q[103],q[102],q[101],q[100],q_b_unconnected_wire_99,q_b_unconnected_wire_98,q_b_unconnected_wire_97,q_b_unconnected_wire_96,q[95],q[94],q[93],q[92],q[91],q[90],q[89],q[88],q[87],q[86],q[85],q[84],q_b_unconnected_wire_83,q_b_unconnected_wire_82,q_b_unconnected_wire_81,q_b_unconnected_wire_80,
q[79],q[78],q[77],q[76],q[75],q[74],q[73],q[72],q[71],q[70],q[69],q[68],q_b_unconnected_wire_67,q_b_unconnected_wire_66,q_b_unconnected_wire_65,q_b_unconnected_wire_64,q[63],q[62],q[61],q[60],q[59],q[58],q[57],q[56],q[55],q[54],q[53],q[52],q_b_unconnected_wire_51,q_b_unconnected_wire_50,q_b_unconnected_wire_49,q_b_unconnected_wire_48,q[47],q[46],q[45],q[44],q[43],q[42],q[41],q[40],q[39],q[38],q[37],q[36],q_b_unconnected_wire_35,
q_b_unconnected_wire_34,q_b_unconnected_wire_33,q_b_unconnected_wire_32,q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,
q_b_unconnected_wire_0}),
	.address_a({\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.clocken1(\valid_rreq~combout ),
	.wren_a(\valid_wreq~combout ),
	.address_b({\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock),
	.data_a({gnd,gnd,data[255],data[254],data[253],data[252],data[251],data[250],data[249],data[248],data[247],data[246],data[245],data[244],gnd,gnd,gnd,gnd,data[239],data[238],data[237],data[236],data[235],data[234],data[233],data[232],data[231],data[230],data[229],data[228],gnd,gnd,gnd,gnd,data[223],data[222],data[221],data[220],data[219],data[218],data[217],data[216],data[215],data[214],data[213],data[212],gnd,gnd,gnd,gnd,data[207],data[206],data[205],data[204],data[203],data[202],data[201],data[200],data[199],data[198],data[197],data[196],gnd,gnd,gnd,gnd,data[191],data[190],
data[189],data[188],data[187],data[186],data[185],data[184],data[183],data[182],data[181],data[180],gnd,gnd,gnd,gnd,data[175],data[174],data[173],data[172],data[171],data[170],data[169],data[168],data[167],data[166],data[165],data[164],gnd,gnd,gnd,gnd,data[159],data[158],data[157],data[156],data[155],data[154],data[153],data[152],data[151],data[150],data[149],data[148],gnd,gnd,gnd,gnd,data[143],data[142],data[141],data[140],data[139],data[138],data[137],data[136],data[135],data[134],data[133],data[132],gnd,gnd,gnd,gnd,data[127],data[126],data[125],data[124],data[123],data[122],
data[121],data[120],data[119],data[118],data[117],data[116],gnd,gnd,gnd,gnd,data[111],data[110],data[109],data[108],data[107],data[106],data[105],data[104],data[103],data[102],data[101],data[100],gnd,gnd,gnd,gnd,data[95],data[94],data[93],data[92],data[91],data[90],data[89],data[88],data[87],data[86],data[85],data[84],gnd,gnd,gnd,gnd,data[79],data[78],data[77],data[76],data[75],data[74],data[73],data[72],data[71],data[70],data[69],data[68],gnd,gnd,gnd,gnd,data[63],data[62],data[61],data[60],data[59],data[58],data[57],data[56],data[55],data[54],
data[53],data[52],gnd,gnd,gnd,gnd,data[47],data[46],data[45],data[44],data[43],data[42],data[41],data[40],data[39],data[38],data[37],data[36],gnd,gnd,gnd,gnd,data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],gnd,gnd,gnd,gnd,data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],gnd,gnd,gnd,gnd}));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\empty_dff~q ),
	.datab(usedw_process),
	.datac(sink_ready_ctrl),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hFEFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb \_~0 (
	.dataa(counter_reg_bit_2),
	.datab(in_valid),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb valid_wreq(
	.dataa(in_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(full_dff1),
	.cin(gnd),
	.combout(\valid_wreq~combout ),
	.cout());
defparam valid_wreq.lut_mask = 16'hAAFF;
defparam valid_wreq.sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hAFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(in_valid),
	.datab(gnd),
	.datac(full_dff1),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hAFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb valid_rreq(
	.dataa(\empty_dff~q ),
	.datab(dffe_nae),
	.datac(sink_ready_ctrl),
	.datad(dffe_af),
	.cin(gnd),
	.combout(\valid_rreq~combout ),
	.cout());
defparam valid_rreq.lut_mask = 16'hFEFF;
defparam valid_rreq.sum_lutc_input = "datac";

cycloneive_lcell_comb \_~1 (
	.dataa(full_dff1),
	.datab(\_~0_combout ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hEEFF;
defparam \_~1 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_1bh1 (
	q_b,
	address_a,
	clocken1,
	wren_a,
	address_b,
	clock1,
	clock0,
	data_a)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q_b;
input 	[2:0] address_a;
input 	clocken1;
input 	wren_a;
input 	[2:0] address_b;
input 	clock1;
input 	clock0;
input 	[257:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a170_PORTBDATAOUT_bus;
wire [143:0] ram_block1a169_PORTBDATAOUT_bus;
wire [143:0] ram_block1a168_PORTBDATAOUT_bus;
wire [143:0] ram_block1a167_PORTBDATAOUT_bus;
wire [143:0] ram_block1a166_PORTBDATAOUT_bus;
wire [143:0] ram_block1a165_PORTBDATAOUT_bus;
wire [143:0] ram_block1a164_PORTBDATAOUT_bus;
wire [143:0] ram_block1a106_PORTBDATAOUT_bus;
wire [143:0] ram_block1a105_PORTBDATAOUT_bus;
wire [143:0] ram_block1a104_PORTBDATAOUT_bus;
wire [143:0] ram_block1a103_PORTBDATAOUT_bus;
wire [143:0] ram_block1a102_PORTBDATAOUT_bus;
wire [143:0] ram_block1a101_PORTBDATAOUT_bus;
wire [143:0] ram_block1a100_PORTBDATAOUT_bus;
wire [143:0] ram_block1a234_PORTBDATAOUT_bus;
wire [143:0] ram_block1a233_PORTBDATAOUT_bus;
wire [143:0] ram_block1a232_PORTBDATAOUT_bus;
wire [143:0] ram_block1a231_PORTBDATAOUT_bus;
wire [143:0] ram_block1a230_PORTBDATAOUT_bus;
wire [143:0] ram_block1a229_PORTBDATAOUT_bus;
wire [143:0] ram_block1a228_PORTBDATAOUT_bus;
wire [143:0] ram_block1a42_PORTBDATAOUT_bus;
wire [143:0] ram_block1a41_PORTBDATAOUT_bus;
wire [143:0] ram_block1a40_PORTBDATAOUT_bus;
wire [143:0] ram_block1a39_PORTBDATAOUT_bus;
wire [143:0] ram_block1a38_PORTBDATAOUT_bus;
wire [143:0] ram_block1a37_PORTBDATAOUT_bus;
wire [143:0] ram_block1a36_PORTBDATAOUT_bus;
wire [143:0] ram_block1a186_PORTBDATAOUT_bus;
wire [143:0] ram_block1a185_PORTBDATAOUT_bus;
wire [143:0] ram_block1a184_PORTBDATAOUT_bus;
wire [143:0] ram_block1a183_PORTBDATAOUT_bus;
wire [143:0] ram_block1a182_PORTBDATAOUT_bus;
wire [143:0] ram_block1a181_PORTBDATAOUT_bus;
wire [143:0] ram_block1a180_PORTBDATAOUT_bus;
wire [143:0] ram_block1a122_PORTBDATAOUT_bus;
wire [143:0] ram_block1a121_PORTBDATAOUT_bus;
wire [143:0] ram_block1a120_PORTBDATAOUT_bus;
wire [143:0] ram_block1a119_PORTBDATAOUT_bus;
wire [143:0] ram_block1a118_PORTBDATAOUT_bus;
wire [143:0] ram_block1a117_PORTBDATAOUT_bus;
wire [143:0] ram_block1a116_PORTBDATAOUT_bus;
wire [143:0] ram_block1a250_PORTBDATAOUT_bus;
wire [143:0] ram_block1a249_PORTBDATAOUT_bus;
wire [143:0] ram_block1a248_PORTBDATAOUT_bus;
wire [143:0] ram_block1a247_PORTBDATAOUT_bus;
wire [143:0] ram_block1a246_PORTBDATAOUT_bus;
wire [143:0] ram_block1a245_PORTBDATAOUT_bus;
wire [143:0] ram_block1a244_PORTBDATAOUT_bus;
wire [143:0] ram_block1a58_PORTBDATAOUT_bus;
wire [143:0] ram_block1a57_PORTBDATAOUT_bus;
wire [143:0] ram_block1a56_PORTBDATAOUT_bus;
wire [143:0] ram_block1a55_PORTBDATAOUT_bus;
wire [143:0] ram_block1a54_PORTBDATAOUT_bus;
wire [143:0] ram_block1a53_PORTBDATAOUT_bus;
wire [143:0] ram_block1a52_PORTBDATAOUT_bus;
wire [143:0] ram_block1a90_PORTBDATAOUT_bus;
wire [143:0] ram_block1a89_PORTBDATAOUT_bus;
wire [143:0] ram_block1a88_PORTBDATAOUT_bus;
wire [143:0] ram_block1a87_PORTBDATAOUT_bus;
wire [143:0] ram_block1a86_PORTBDATAOUT_bus;
wire [143:0] ram_block1a85_PORTBDATAOUT_bus;
wire [143:0] ram_block1a84_PORTBDATAOUT_bus;
wire [143:0] ram_block1a154_PORTBDATAOUT_bus;
wire [143:0] ram_block1a153_PORTBDATAOUT_bus;
wire [143:0] ram_block1a152_PORTBDATAOUT_bus;
wire [143:0] ram_block1a151_PORTBDATAOUT_bus;
wire [143:0] ram_block1a150_PORTBDATAOUT_bus;
wire [143:0] ram_block1a149_PORTBDATAOUT_bus;
wire [143:0] ram_block1a148_PORTBDATAOUT_bus;
wire [143:0] ram_block1a218_PORTBDATAOUT_bus;
wire [143:0] ram_block1a217_PORTBDATAOUT_bus;
wire [143:0] ram_block1a216_PORTBDATAOUT_bus;
wire [143:0] ram_block1a215_PORTBDATAOUT_bus;
wire [143:0] ram_block1a214_PORTBDATAOUT_bus;
wire [143:0] ram_block1a213_PORTBDATAOUT_bus;
wire [143:0] ram_block1a212_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a74_PORTBDATAOUT_bus;
wire [143:0] ram_block1a73_PORTBDATAOUT_bus;
wire [143:0] ram_block1a72_PORTBDATAOUT_bus;
wire [143:0] ram_block1a71_PORTBDATAOUT_bus;
wire [143:0] ram_block1a70_PORTBDATAOUT_bus;
wire [143:0] ram_block1a69_PORTBDATAOUT_bus;
wire [143:0] ram_block1a68_PORTBDATAOUT_bus;
wire [143:0] ram_block1a138_PORTBDATAOUT_bus;
wire [143:0] ram_block1a137_PORTBDATAOUT_bus;
wire [143:0] ram_block1a136_PORTBDATAOUT_bus;
wire [143:0] ram_block1a135_PORTBDATAOUT_bus;
wire [143:0] ram_block1a134_PORTBDATAOUT_bus;
wire [143:0] ram_block1a133_PORTBDATAOUT_bus;
wire [143:0] ram_block1a132_PORTBDATAOUT_bus;
wire [143:0] ram_block1a202_PORTBDATAOUT_bus;
wire [143:0] ram_block1a201_PORTBDATAOUT_bus;
wire [143:0] ram_block1a200_PORTBDATAOUT_bus;
wire [143:0] ram_block1a199_PORTBDATAOUT_bus;
wire [143:0] ram_block1a198_PORTBDATAOUT_bus;
wire [143:0] ram_block1a197_PORTBDATAOUT_bus;
wire [143:0] ram_block1a196_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a107_PORTBDATAOUT_bus;
wire [143:0] ram_block1a123_PORTBDATAOUT_bus;
wire [143:0] ram_block1a91_PORTBDATAOUT_bus;
wire [143:0] ram_block1a75_PORTBDATAOUT_bus;
wire [143:0] ram_block1a171_PORTBDATAOUT_bus;
wire [143:0] ram_block1a187_PORTBDATAOUT_bus;
wire [143:0] ram_block1a155_PORTBDATAOUT_bus;
wire [143:0] ram_block1a139_PORTBDATAOUT_bus;
wire [143:0] ram_block1a235_PORTBDATAOUT_bus;
wire [143:0] ram_block1a251_PORTBDATAOUT_bus;
wire [143:0] ram_block1a219_PORTBDATAOUT_bus;
wire [143:0] ram_block1a203_PORTBDATAOUT_bus;
wire [143:0] ram_block1a43_PORTBDATAOUT_bus;
wire [143:0] ram_block1a59_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a108_PORTBDATAOUT_bus;
wire [143:0] ram_block1a172_PORTBDATAOUT_bus;
wire [143:0] ram_block1a236_PORTBDATAOUT_bus;
wire [143:0] ram_block1a44_PORTBDATAOUT_bus;
wire [143:0] ram_block1a124_PORTBDATAOUT_bus;
wire [143:0] ram_block1a188_PORTBDATAOUT_bus;
wire [143:0] ram_block1a252_PORTBDATAOUT_bus;
wire [143:0] ram_block1a60_PORTBDATAOUT_bus;
wire [143:0] ram_block1a156_PORTBDATAOUT_bus;
wire [143:0] ram_block1a92_PORTBDATAOUT_bus;
wire [143:0] ram_block1a220_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a140_PORTBDATAOUT_bus;
wire [143:0] ram_block1a76_PORTBDATAOUT_bus;
wire [143:0] ram_block1a204_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a173_PORTBDATAOUT_bus;
wire [143:0] ram_block1a189_PORTBDATAOUT_bus;
wire [143:0] ram_block1a157_PORTBDATAOUT_bus;
wire [143:0] ram_block1a141_PORTBDATAOUT_bus;
wire [143:0] ram_block1a109_PORTBDATAOUT_bus;
wire [143:0] ram_block1a125_PORTBDATAOUT_bus;
wire [143:0] ram_block1a93_PORTBDATAOUT_bus;
wire [143:0] ram_block1a77_PORTBDATAOUT_bus;
wire [143:0] ram_block1a237_PORTBDATAOUT_bus;
wire [143:0] ram_block1a253_PORTBDATAOUT_bus;
wire [143:0] ram_block1a221_PORTBDATAOUT_bus;
wire [143:0] ram_block1a205_PORTBDATAOUT_bus;
wire [143:0] ram_block1a45_PORTBDATAOUT_bus;
wire [143:0] ram_block1a61_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a174_PORTBDATAOUT_bus;
wire [143:0] ram_block1a110_PORTBDATAOUT_bus;
wire [143:0] ram_block1a238_PORTBDATAOUT_bus;
wire [143:0] ram_block1a46_PORTBDATAOUT_bus;
wire [143:0] ram_block1a190_PORTBDATAOUT_bus;
wire [143:0] ram_block1a126_PORTBDATAOUT_bus;
wire [143:0] ram_block1a254_PORTBDATAOUT_bus;
wire [143:0] ram_block1a62_PORTBDATAOUT_bus;
wire [143:0] ram_block1a94_PORTBDATAOUT_bus;
wire [143:0] ram_block1a158_PORTBDATAOUT_bus;
wire [143:0] ram_block1a222_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a78_PORTBDATAOUT_bus;
wire [143:0] ram_block1a142_PORTBDATAOUT_bus;
wire [143:0] ram_block1a206_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a111_PORTBDATAOUT_bus;
wire [143:0] ram_block1a127_PORTBDATAOUT_bus;
wire [143:0] ram_block1a95_PORTBDATAOUT_bus;
wire [143:0] ram_block1a79_PORTBDATAOUT_bus;
wire [143:0] ram_block1a175_PORTBDATAOUT_bus;
wire [143:0] ram_block1a191_PORTBDATAOUT_bus;
wire [143:0] ram_block1a159_PORTBDATAOUT_bus;
wire [143:0] ram_block1a143_PORTBDATAOUT_bus;
wire [143:0] ram_block1a239_PORTBDATAOUT_bus;
wire [143:0] ram_block1a255_PORTBDATAOUT_bus;
wire [143:0] ram_block1a223_PORTBDATAOUT_bus;
wire [143:0] ram_block1a207_PORTBDATAOUT_bus;
wire [143:0] ram_block1a47_PORTBDATAOUT_bus;
wire [143:0] ram_block1a63_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;

assign q_b[170] = ram_block1a170_PORTBDATAOUT_bus[0];

assign q_b[169] = ram_block1a169_PORTBDATAOUT_bus[0];

assign q_b[168] = ram_block1a168_PORTBDATAOUT_bus[0];

assign q_b[167] = ram_block1a167_PORTBDATAOUT_bus[0];

assign q_b[166] = ram_block1a166_PORTBDATAOUT_bus[0];

assign q_b[165] = ram_block1a165_PORTBDATAOUT_bus[0];

assign q_b[164] = ram_block1a164_PORTBDATAOUT_bus[0];

assign q_b[106] = ram_block1a106_PORTBDATAOUT_bus[0];

assign q_b[105] = ram_block1a105_PORTBDATAOUT_bus[0];

assign q_b[104] = ram_block1a104_PORTBDATAOUT_bus[0];

assign q_b[103] = ram_block1a103_PORTBDATAOUT_bus[0];

assign q_b[102] = ram_block1a102_PORTBDATAOUT_bus[0];

assign q_b[101] = ram_block1a101_PORTBDATAOUT_bus[0];

assign q_b[100] = ram_block1a100_PORTBDATAOUT_bus[0];

assign q_b[234] = ram_block1a234_PORTBDATAOUT_bus[0];

assign q_b[233] = ram_block1a233_PORTBDATAOUT_bus[0];

assign q_b[232] = ram_block1a232_PORTBDATAOUT_bus[0];

assign q_b[231] = ram_block1a231_PORTBDATAOUT_bus[0];

assign q_b[230] = ram_block1a230_PORTBDATAOUT_bus[0];

assign q_b[229] = ram_block1a229_PORTBDATAOUT_bus[0];

assign q_b[228] = ram_block1a228_PORTBDATAOUT_bus[0];

assign q_b[42] = ram_block1a42_PORTBDATAOUT_bus[0];

assign q_b[41] = ram_block1a41_PORTBDATAOUT_bus[0];

assign q_b[40] = ram_block1a40_PORTBDATAOUT_bus[0];

assign q_b[39] = ram_block1a39_PORTBDATAOUT_bus[0];

assign q_b[38] = ram_block1a38_PORTBDATAOUT_bus[0];

assign q_b[37] = ram_block1a37_PORTBDATAOUT_bus[0];

assign q_b[36] = ram_block1a36_PORTBDATAOUT_bus[0];

assign q_b[186] = ram_block1a186_PORTBDATAOUT_bus[0];

assign q_b[185] = ram_block1a185_PORTBDATAOUT_bus[0];

assign q_b[184] = ram_block1a184_PORTBDATAOUT_bus[0];

assign q_b[183] = ram_block1a183_PORTBDATAOUT_bus[0];

assign q_b[182] = ram_block1a182_PORTBDATAOUT_bus[0];

assign q_b[181] = ram_block1a181_PORTBDATAOUT_bus[0];

assign q_b[180] = ram_block1a180_PORTBDATAOUT_bus[0];

assign q_b[122] = ram_block1a122_PORTBDATAOUT_bus[0];

assign q_b[121] = ram_block1a121_PORTBDATAOUT_bus[0];

assign q_b[120] = ram_block1a120_PORTBDATAOUT_bus[0];

assign q_b[119] = ram_block1a119_PORTBDATAOUT_bus[0];

assign q_b[118] = ram_block1a118_PORTBDATAOUT_bus[0];

assign q_b[117] = ram_block1a117_PORTBDATAOUT_bus[0];

assign q_b[116] = ram_block1a116_PORTBDATAOUT_bus[0];

assign q_b[250] = ram_block1a250_PORTBDATAOUT_bus[0];

assign q_b[249] = ram_block1a249_PORTBDATAOUT_bus[0];

assign q_b[248] = ram_block1a248_PORTBDATAOUT_bus[0];

assign q_b[247] = ram_block1a247_PORTBDATAOUT_bus[0];

assign q_b[246] = ram_block1a246_PORTBDATAOUT_bus[0];

assign q_b[245] = ram_block1a245_PORTBDATAOUT_bus[0];

assign q_b[244] = ram_block1a244_PORTBDATAOUT_bus[0];

assign q_b[58] = ram_block1a58_PORTBDATAOUT_bus[0];

assign q_b[57] = ram_block1a57_PORTBDATAOUT_bus[0];

assign q_b[56] = ram_block1a56_PORTBDATAOUT_bus[0];

assign q_b[55] = ram_block1a55_PORTBDATAOUT_bus[0];

assign q_b[54] = ram_block1a54_PORTBDATAOUT_bus[0];

assign q_b[53] = ram_block1a53_PORTBDATAOUT_bus[0];

assign q_b[52] = ram_block1a52_PORTBDATAOUT_bus[0];

assign q_b[90] = ram_block1a90_PORTBDATAOUT_bus[0];

assign q_b[89] = ram_block1a89_PORTBDATAOUT_bus[0];

assign q_b[88] = ram_block1a88_PORTBDATAOUT_bus[0];

assign q_b[87] = ram_block1a87_PORTBDATAOUT_bus[0];

assign q_b[86] = ram_block1a86_PORTBDATAOUT_bus[0];

assign q_b[85] = ram_block1a85_PORTBDATAOUT_bus[0];

assign q_b[84] = ram_block1a84_PORTBDATAOUT_bus[0];

assign q_b[154] = ram_block1a154_PORTBDATAOUT_bus[0];

assign q_b[153] = ram_block1a153_PORTBDATAOUT_bus[0];

assign q_b[152] = ram_block1a152_PORTBDATAOUT_bus[0];

assign q_b[151] = ram_block1a151_PORTBDATAOUT_bus[0];

assign q_b[150] = ram_block1a150_PORTBDATAOUT_bus[0];

assign q_b[149] = ram_block1a149_PORTBDATAOUT_bus[0];

assign q_b[148] = ram_block1a148_PORTBDATAOUT_bus[0];

assign q_b[218] = ram_block1a218_PORTBDATAOUT_bus[0];

assign q_b[217] = ram_block1a217_PORTBDATAOUT_bus[0];

assign q_b[216] = ram_block1a216_PORTBDATAOUT_bus[0];

assign q_b[215] = ram_block1a215_PORTBDATAOUT_bus[0];

assign q_b[214] = ram_block1a214_PORTBDATAOUT_bus[0];

assign q_b[213] = ram_block1a213_PORTBDATAOUT_bus[0];

assign q_b[212] = ram_block1a212_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[74] = ram_block1a74_PORTBDATAOUT_bus[0];

assign q_b[73] = ram_block1a73_PORTBDATAOUT_bus[0];

assign q_b[72] = ram_block1a72_PORTBDATAOUT_bus[0];

assign q_b[71] = ram_block1a71_PORTBDATAOUT_bus[0];

assign q_b[70] = ram_block1a70_PORTBDATAOUT_bus[0];

assign q_b[69] = ram_block1a69_PORTBDATAOUT_bus[0];

assign q_b[68] = ram_block1a68_PORTBDATAOUT_bus[0];

assign q_b[138] = ram_block1a138_PORTBDATAOUT_bus[0];

assign q_b[137] = ram_block1a137_PORTBDATAOUT_bus[0];

assign q_b[136] = ram_block1a136_PORTBDATAOUT_bus[0];

assign q_b[135] = ram_block1a135_PORTBDATAOUT_bus[0];

assign q_b[134] = ram_block1a134_PORTBDATAOUT_bus[0];

assign q_b[133] = ram_block1a133_PORTBDATAOUT_bus[0];

assign q_b[132] = ram_block1a132_PORTBDATAOUT_bus[0];

assign q_b[202] = ram_block1a202_PORTBDATAOUT_bus[0];

assign q_b[201] = ram_block1a201_PORTBDATAOUT_bus[0];

assign q_b[200] = ram_block1a200_PORTBDATAOUT_bus[0];

assign q_b[199] = ram_block1a199_PORTBDATAOUT_bus[0];

assign q_b[198] = ram_block1a198_PORTBDATAOUT_bus[0];

assign q_b[197] = ram_block1a197_PORTBDATAOUT_bus[0];

assign q_b[196] = ram_block1a196_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[107] = ram_block1a107_PORTBDATAOUT_bus[0];

assign q_b[123] = ram_block1a123_PORTBDATAOUT_bus[0];

assign q_b[91] = ram_block1a91_PORTBDATAOUT_bus[0];

assign q_b[75] = ram_block1a75_PORTBDATAOUT_bus[0];

assign q_b[171] = ram_block1a171_PORTBDATAOUT_bus[0];

assign q_b[187] = ram_block1a187_PORTBDATAOUT_bus[0];

assign q_b[155] = ram_block1a155_PORTBDATAOUT_bus[0];

assign q_b[139] = ram_block1a139_PORTBDATAOUT_bus[0];

assign q_b[235] = ram_block1a235_PORTBDATAOUT_bus[0];

assign q_b[251] = ram_block1a251_PORTBDATAOUT_bus[0];

assign q_b[219] = ram_block1a219_PORTBDATAOUT_bus[0];

assign q_b[203] = ram_block1a203_PORTBDATAOUT_bus[0];

assign q_b[43] = ram_block1a43_PORTBDATAOUT_bus[0];

assign q_b[59] = ram_block1a59_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[108] = ram_block1a108_PORTBDATAOUT_bus[0];

assign q_b[172] = ram_block1a172_PORTBDATAOUT_bus[0];

assign q_b[236] = ram_block1a236_PORTBDATAOUT_bus[0];

assign q_b[44] = ram_block1a44_PORTBDATAOUT_bus[0];

assign q_b[124] = ram_block1a124_PORTBDATAOUT_bus[0];

assign q_b[188] = ram_block1a188_PORTBDATAOUT_bus[0];

assign q_b[252] = ram_block1a252_PORTBDATAOUT_bus[0];

assign q_b[60] = ram_block1a60_PORTBDATAOUT_bus[0];

assign q_b[156] = ram_block1a156_PORTBDATAOUT_bus[0];

assign q_b[92] = ram_block1a92_PORTBDATAOUT_bus[0];

assign q_b[220] = ram_block1a220_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[140] = ram_block1a140_PORTBDATAOUT_bus[0];

assign q_b[76] = ram_block1a76_PORTBDATAOUT_bus[0];

assign q_b[204] = ram_block1a204_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[173] = ram_block1a173_PORTBDATAOUT_bus[0];

assign q_b[189] = ram_block1a189_PORTBDATAOUT_bus[0];

assign q_b[157] = ram_block1a157_PORTBDATAOUT_bus[0];

assign q_b[141] = ram_block1a141_PORTBDATAOUT_bus[0];

assign q_b[109] = ram_block1a109_PORTBDATAOUT_bus[0];

assign q_b[125] = ram_block1a125_PORTBDATAOUT_bus[0];

assign q_b[93] = ram_block1a93_PORTBDATAOUT_bus[0];

assign q_b[77] = ram_block1a77_PORTBDATAOUT_bus[0];

assign q_b[237] = ram_block1a237_PORTBDATAOUT_bus[0];

assign q_b[253] = ram_block1a253_PORTBDATAOUT_bus[0];

assign q_b[221] = ram_block1a221_PORTBDATAOUT_bus[0];

assign q_b[205] = ram_block1a205_PORTBDATAOUT_bus[0];

assign q_b[45] = ram_block1a45_PORTBDATAOUT_bus[0];

assign q_b[61] = ram_block1a61_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[174] = ram_block1a174_PORTBDATAOUT_bus[0];

assign q_b[110] = ram_block1a110_PORTBDATAOUT_bus[0];

assign q_b[238] = ram_block1a238_PORTBDATAOUT_bus[0];

assign q_b[46] = ram_block1a46_PORTBDATAOUT_bus[0];

assign q_b[190] = ram_block1a190_PORTBDATAOUT_bus[0];

assign q_b[126] = ram_block1a126_PORTBDATAOUT_bus[0];

assign q_b[254] = ram_block1a254_PORTBDATAOUT_bus[0];

assign q_b[62] = ram_block1a62_PORTBDATAOUT_bus[0];

assign q_b[94] = ram_block1a94_PORTBDATAOUT_bus[0];

assign q_b[158] = ram_block1a158_PORTBDATAOUT_bus[0];

assign q_b[222] = ram_block1a222_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[78] = ram_block1a78_PORTBDATAOUT_bus[0];

assign q_b[142] = ram_block1a142_PORTBDATAOUT_bus[0];

assign q_b[206] = ram_block1a206_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[111] = ram_block1a111_PORTBDATAOUT_bus[0];

assign q_b[127] = ram_block1a127_PORTBDATAOUT_bus[0];

assign q_b[95] = ram_block1a95_PORTBDATAOUT_bus[0];

assign q_b[79] = ram_block1a79_PORTBDATAOUT_bus[0];

assign q_b[175] = ram_block1a175_PORTBDATAOUT_bus[0];

assign q_b[191] = ram_block1a191_PORTBDATAOUT_bus[0];

assign q_b[159] = ram_block1a159_PORTBDATAOUT_bus[0];

assign q_b[143] = ram_block1a143_PORTBDATAOUT_bus[0];

assign q_b[239] = ram_block1a239_PORTBDATAOUT_bus[0];

assign q_b[255] = ram_block1a255_PORTBDATAOUT_bus[0];

assign q_b[223] = ram_block1a223_PORTBDATAOUT_bus[0];

assign q_b[207] = ram_block1a207_PORTBDATAOUT_bus[0];

assign q_b[47] = ram_block1a47_PORTBDATAOUT_bus[0];

assign q_b[63] = ram_block1a63_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a170(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[170]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a170_PORTBDATAOUT_bus));
defparam ram_block1a170.clk1_output_clock_enable = "ena1";
defparam ram_block1a170.data_interleave_offset_in_bits = 1;
defparam ram_block1a170.data_interleave_width_in_bits = 1;
defparam ram_block1a170.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a170.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a170.operation_mode = "dual_port";
defparam ram_block1a170.port_a_address_clear = "none";
defparam ram_block1a170.port_a_address_width = 3;
defparam ram_block1a170.port_a_data_out_clear = "none";
defparam ram_block1a170.port_a_data_out_clock = "none";
defparam ram_block1a170.port_a_data_width = 1;
defparam ram_block1a170.port_a_first_address = 0;
defparam ram_block1a170.port_a_first_bit_number = 170;
defparam ram_block1a170.port_a_last_address = 7;
defparam ram_block1a170.port_a_logical_ram_depth = 8;
defparam ram_block1a170.port_a_logical_ram_width = 258;
defparam ram_block1a170.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a170.port_b_address_clear = "none";
defparam ram_block1a170.port_b_address_clock = "clock1";
defparam ram_block1a170.port_b_address_width = 3;
defparam ram_block1a170.port_b_data_out_clear = "none";
defparam ram_block1a170.port_b_data_out_clock = "clock1";
defparam ram_block1a170.port_b_data_width = 1;
defparam ram_block1a170.port_b_first_address = 0;
defparam ram_block1a170.port_b_first_bit_number = 170;
defparam ram_block1a170.port_b_last_address = 7;
defparam ram_block1a170.port_b_logical_ram_depth = 8;
defparam ram_block1a170.port_b_logical_ram_width = 258;
defparam ram_block1a170.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a170.port_b_read_enable_clock = "clock1";
defparam ram_block1a170.ram_block_type = "auto";

cycloneive_ram_block ram_block1a169(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[169]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a169_PORTBDATAOUT_bus));
defparam ram_block1a169.clk1_output_clock_enable = "ena1";
defparam ram_block1a169.data_interleave_offset_in_bits = 1;
defparam ram_block1a169.data_interleave_width_in_bits = 1;
defparam ram_block1a169.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a169.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a169.operation_mode = "dual_port";
defparam ram_block1a169.port_a_address_clear = "none";
defparam ram_block1a169.port_a_address_width = 3;
defparam ram_block1a169.port_a_data_out_clear = "none";
defparam ram_block1a169.port_a_data_out_clock = "none";
defparam ram_block1a169.port_a_data_width = 1;
defparam ram_block1a169.port_a_first_address = 0;
defparam ram_block1a169.port_a_first_bit_number = 169;
defparam ram_block1a169.port_a_last_address = 7;
defparam ram_block1a169.port_a_logical_ram_depth = 8;
defparam ram_block1a169.port_a_logical_ram_width = 258;
defparam ram_block1a169.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a169.port_b_address_clear = "none";
defparam ram_block1a169.port_b_address_clock = "clock1";
defparam ram_block1a169.port_b_address_width = 3;
defparam ram_block1a169.port_b_data_out_clear = "none";
defparam ram_block1a169.port_b_data_out_clock = "clock1";
defparam ram_block1a169.port_b_data_width = 1;
defparam ram_block1a169.port_b_first_address = 0;
defparam ram_block1a169.port_b_first_bit_number = 169;
defparam ram_block1a169.port_b_last_address = 7;
defparam ram_block1a169.port_b_logical_ram_depth = 8;
defparam ram_block1a169.port_b_logical_ram_width = 258;
defparam ram_block1a169.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a169.port_b_read_enable_clock = "clock1";
defparam ram_block1a169.ram_block_type = "auto";

cycloneive_ram_block ram_block1a168(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[168]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a168_PORTBDATAOUT_bus));
defparam ram_block1a168.clk1_output_clock_enable = "ena1";
defparam ram_block1a168.data_interleave_offset_in_bits = 1;
defparam ram_block1a168.data_interleave_width_in_bits = 1;
defparam ram_block1a168.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a168.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a168.operation_mode = "dual_port";
defparam ram_block1a168.port_a_address_clear = "none";
defparam ram_block1a168.port_a_address_width = 3;
defparam ram_block1a168.port_a_data_out_clear = "none";
defparam ram_block1a168.port_a_data_out_clock = "none";
defparam ram_block1a168.port_a_data_width = 1;
defparam ram_block1a168.port_a_first_address = 0;
defparam ram_block1a168.port_a_first_bit_number = 168;
defparam ram_block1a168.port_a_last_address = 7;
defparam ram_block1a168.port_a_logical_ram_depth = 8;
defparam ram_block1a168.port_a_logical_ram_width = 258;
defparam ram_block1a168.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a168.port_b_address_clear = "none";
defparam ram_block1a168.port_b_address_clock = "clock1";
defparam ram_block1a168.port_b_address_width = 3;
defparam ram_block1a168.port_b_data_out_clear = "none";
defparam ram_block1a168.port_b_data_out_clock = "clock1";
defparam ram_block1a168.port_b_data_width = 1;
defparam ram_block1a168.port_b_first_address = 0;
defparam ram_block1a168.port_b_first_bit_number = 168;
defparam ram_block1a168.port_b_last_address = 7;
defparam ram_block1a168.port_b_logical_ram_depth = 8;
defparam ram_block1a168.port_b_logical_ram_width = 258;
defparam ram_block1a168.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a168.port_b_read_enable_clock = "clock1";
defparam ram_block1a168.ram_block_type = "auto";

cycloneive_ram_block ram_block1a167(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[167]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a167_PORTBDATAOUT_bus));
defparam ram_block1a167.clk1_output_clock_enable = "ena1";
defparam ram_block1a167.data_interleave_offset_in_bits = 1;
defparam ram_block1a167.data_interleave_width_in_bits = 1;
defparam ram_block1a167.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a167.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a167.operation_mode = "dual_port";
defparam ram_block1a167.port_a_address_clear = "none";
defparam ram_block1a167.port_a_address_width = 3;
defparam ram_block1a167.port_a_data_out_clear = "none";
defparam ram_block1a167.port_a_data_out_clock = "none";
defparam ram_block1a167.port_a_data_width = 1;
defparam ram_block1a167.port_a_first_address = 0;
defparam ram_block1a167.port_a_first_bit_number = 167;
defparam ram_block1a167.port_a_last_address = 7;
defparam ram_block1a167.port_a_logical_ram_depth = 8;
defparam ram_block1a167.port_a_logical_ram_width = 258;
defparam ram_block1a167.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a167.port_b_address_clear = "none";
defparam ram_block1a167.port_b_address_clock = "clock1";
defparam ram_block1a167.port_b_address_width = 3;
defparam ram_block1a167.port_b_data_out_clear = "none";
defparam ram_block1a167.port_b_data_out_clock = "clock1";
defparam ram_block1a167.port_b_data_width = 1;
defparam ram_block1a167.port_b_first_address = 0;
defparam ram_block1a167.port_b_first_bit_number = 167;
defparam ram_block1a167.port_b_last_address = 7;
defparam ram_block1a167.port_b_logical_ram_depth = 8;
defparam ram_block1a167.port_b_logical_ram_width = 258;
defparam ram_block1a167.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a167.port_b_read_enable_clock = "clock1";
defparam ram_block1a167.ram_block_type = "auto";

cycloneive_ram_block ram_block1a166(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[166]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a166_PORTBDATAOUT_bus));
defparam ram_block1a166.clk1_output_clock_enable = "ena1";
defparam ram_block1a166.data_interleave_offset_in_bits = 1;
defparam ram_block1a166.data_interleave_width_in_bits = 1;
defparam ram_block1a166.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a166.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a166.operation_mode = "dual_port";
defparam ram_block1a166.port_a_address_clear = "none";
defparam ram_block1a166.port_a_address_width = 3;
defparam ram_block1a166.port_a_data_out_clear = "none";
defparam ram_block1a166.port_a_data_out_clock = "none";
defparam ram_block1a166.port_a_data_width = 1;
defparam ram_block1a166.port_a_first_address = 0;
defparam ram_block1a166.port_a_first_bit_number = 166;
defparam ram_block1a166.port_a_last_address = 7;
defparam ram_block1a166.port_a_logical_ram_depth = 8;
defparam ram_block1a166.port_a_logical_ram_width = 258;
defparam ram_block1a166.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a166.port_b_address_clear = "none";
defparam ram_block1a166.port_b_address_clock = "clock1";
defparam ram_block1a166.port_b_address_width = 3;
defparam ram_block1a166.port_b_data_out_clear = "none";
defparam ram_block1a166.port_b_data_out_clock = "clock1";
defparam ram_block1a166.port_b_data_width = 1;
defparam ram_block1a166.port_b_first_address = 0;
defparam ram_block1a166.port_b_first_bit_number = 166;
defparam ram_block1a166.port_b_last_address = 7;
defparam ram_block1a166.port_b_logical_ram_depth = 8;
defparam ram_block1a166.port_b_logical_ram_width = 258;
defparam ram_block1a166.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a166.port_b_read_enable_clock = "clock1";
defparam ram_block1a166.ram_block_type = "auto";

cycloneive_ram_block ram_block1a165(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[165]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a165_PORTBDATAOUT_bus));
defparam ram_block1a165.clk1_output_clock_enable = "ena1";
defparam ram_block1a165.data_interleave_offset_in_bits = 1;
defparam ram_block1a165.data_interleave_width_in_bits = 1;
defparam ram_block1a165.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a165.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a165.operation_mode = "dual_port";
defparam ram_block1a165.port_a_address_clear = "none";
defparam ram_block1a165.port_a_address_width = 3;
defparam ram_block1a165.port_a_data_out_clear = "none";
defparam ram_block1a165.port_a_data_out_clock = "none";
defparam ram_block1a165.port_a_data_width = 1;
defparam ram_block1a165.port_a_first_address = 0;
defparam ram_block1a165.port_a_first_bit_number = 165;
defparam ram_block1a165.port_a_last_address = 7;
defparam ram_block1a165.port_a_logical_ram_depth = 8;
defparam ram_block1a165.port_a_logical_ram_width = 258;
defparam ram_block1a165.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a165.port_b_address_clear = "none";
defparam ram_block1a165.port_b_address_clock = "clock1";
defparam ram_block1a165.port_b_address_width = 3;
defparam ram_block1a165.port_b_data_out_clear = "none";
defparam ram_block1a165.port_b_data_out_clock = "clock1";
defparam ram_block1a165.port_b_data_width = 1;
defparam ram_block1a165.port_b_first_address = 0;
defparam ram_block1a165.port_b_first_bit_number = 165;
defparam ram_block1a165.port_b_last_address = 7;
defparam ram_block1a165.port_b_logical_ram_depth = 8;
defparam ram_block1a165.port_b_logical_ram_width = 258;
defparam ram_block1a165.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a165.port_b_read_enable_clock = "clock1";
defparam ram_block1a165.ram_block_type = "auto";

cycloneive_ram_block ram_block1a164(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[164]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a164_PORTBDATAOUT_bus));
defparam ram_block1a164.clk1_output_clock_enable = "ena1";
defparam ram_block1a164.data_interleave_offset_in_bits = 1;
defparam ram_block1a164.data_interleave_width_in_bits = 1;
defparam ram_block1a164.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a164.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a164.operation_mode = "dual_port";
defparam ram_block1a164.port_a_address_clear = "none";
defparam ram_block1a164.port_a_address_width = 3;
defparam ram_block1a164.port_a_data_out_clear = "none";
defparam ram_block1a164.port_a_data_out_clock = "none";
defparam ram_block1a164.port_a_data_width = 1;
defparam ram_block1a164.port_a_first_address = 0;
defparam ram_block1a164.port_a_first_bit_number = 164;
defparam ram_block1a164.port_a_last_address = 7;
defparam ram_block1a164.port_a_logical_ram_depth = 8;
defparam ram_block1a164.port_a_logical_ram_width = 258;
defparam ram_block1a164.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a164.port_b_address_clear = "none";
defparam ram_block1a164.port_b_address_clock = "clock1";
defparam ram_block1a164.port_b_address_width = 3;
defparam ram_block1a164.port_b_data_out_clear = "none";
defparam ram_block1a164.port_b_data_out_clock = "clock1";
defparam ram_block1a164.port_b_data_width = 1;
defparam ram_block1a164.port_b_first_address = 0;
defparam ram_block1a164.port_b_first_bit_number = 164;
defparam ram_block1a164.port_b_last_address = 7;
defparam ram_block1a164.port_b_logical_ram_depth = 8;
defparam ram_block1a164.port_b_logical_ram_width = 258;
defparam ram_block1a164.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a164.port_b_read_enable_clock = "clock1";
defparam ram_block1a164.ram_block_type = "auto";

cycloneive_ram_block ram_block1a106(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[106]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a106_PORTBDATAOUT_bus));
defparam ram_block1a106.clk1_output_clock_enable = "ena1";
defparam ram_block1a106.data_interleave_offset_in_bits = 1;
defparam ram_block1a106.data_interleave_width_in_bits = 1;
defparam ram_block1a106.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a106.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a106.operation_mode = "dual_port";
defparam ram_block1a106.port_a_address_clear = "none";
defparam ram_block1a106.port_a_address_width = 3;
defparam ram_block1a106.port_a_data_out_clear = "none";
defparam ram_block1a106.port_a_data_out_clock = "none";
defparam ram_block1a106.port_a_data_width = 1;
defparam ram_block1a106.port_a_first_address = 0;
defparam ram_block1a106.port_a_first_bit_number = 106;
defparam ram_block1a106.port_a_last_address = 7;
defparam ram_block1a106.port_a_logical_ram_depth = 8;
defparam ram_block1a106.port_a_logical_ram_width = 258;
defparam ram_block1a106.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a106.port_b_address_clear = "none";
defparam ram_block1a106.port_b_address_clock = "clock1";
defparam ram_block1a106.port_b_address_width = 3;
defparam ram_block1a106.port_b_data_out_clear = "none";
defparam ram_block1a106.port_b_data_out_clock = "clock1";
defparam ram_block1a106.port_b_data_width = 1;
defparam ram_block1a106.port_b_first_address = 0;
defparam ram_block1a106.port_b_first_bit_number = 106;
defparam ram_block1a106.port_b_last_address = 7;
defparam ram_block1a106.port_b_logical_ram_depth = 8;
defparam ram_block1a106.port_b_logical_ram_width = 258;
defparam ram_block1a106.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a106.port_b_read_enable_clock = "clock1";
defparam ram_block1a106.ram_block_type = "auto";

cycloneive_ram_block ram_block1a105(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[105]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a105_PORTBDATAOUT_bus));
defparam ram_block1a105.clk1_output_clock_enable = "ena1";
defparam ram_block1a105.data_interleave_offset_in_bits = 1;
defparam ram_block1a105.data_interleave_width_in_bits = 1;
defparam ram_block1a105.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a105.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a105.operation_mode = "dual_port";
defparam ram_block1a105.port_a_address_clear = "none";
defparam ram_block1a105.port_a_address_width = 3;
defparam ram_block1a105.port_a_data_out_clear = "none";
defparam ram_block1a105.port_a_data_out_clock = "none";
defparam ram_block1a105.port_a_data_width = 1;
defparam ram_block1a105.port_a_first_address = 0;
defparam ram_block1a105.port_a_first_bit_number = 105;
defparam ram_block1a105.port_a_last_address = 7;
defparam ram_block1a105.port_a_logical_ram_depth = 8;
defparam ram_block1a105.port_a_logical_ram_width = 258;
defparam ram_block1a105.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a105.port_b_address_clear = "none";
defparam ram_block1a105.port_b_address_clock = "clock1";
defparam ram_block1a105.port_b_address_width = 3;
defparam ram_block1a105.port_b_data_out_clear = "none";
defparam ram_block1a105.port_b_data_out_clock = "clock1";
defparam ram_block1a105.port_b_data_width = 1;
defparam ram_block1a105.port_b_first_address = 0;
defparam ram_block1a105.port_b_first_bit_number = 105;
defparam ram_block1a105.port_b_last_address = 7;
defparam ram_block1a105.port_b_logical_ram_depth = 8;
defparam ram_block1a105.port_b_logical_ram_width = 258;
defparam ram_block1a105.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a105.port_b_read_enable_clock = "clock1";
defparam ram_block1a105.ram_block_type = "auto";

cycloneive_ram_block ram_block1a104(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[104]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a104_PORTBDATAOUT_bus));
defparam ram_block1a104.clk1_output_clock_enable = "ena1";
defparam ram_block1a104.data_interleave_offset_in_bits = 1;
defparam ram_block1a104.data_interleave_width_in_bits = 1;
defparam ram_block1a104.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a104.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a104.operation_mode = "dual_port";
defparam ram_block1a104.port_a_address_clear = "none";
defparam ram_block1a104.port_a_address_width = 3;
defparam ram_block1a104.port_a_data_out_clear = "none";
defparam ram_block1a104.port_a_data_out_clock = "none";
defparam ram_block1a104.port_a_data_width = 1;
defparam ram_block1a104.port_a_first_address = 0;
defparam ram_block1a104.port_a_first_bit_number = 104;
defparam ram_block1a104.port_a_last_address = 7;
defparam ram_block1a104.port_a_logical_ram_depth = 8;
defparam ram_block1a104.port_a_logical_ram_width = 258;
defparam ram_block1a104.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a104.port_b_address_clear = "none";
defparam ram_block1a104.port_b_address_clock = "clock1";
defparam ram_block1a104.port_b_address_width = 3;
defparam ram_block1a104.port_b_data_out_clear = "none";
defparam ram_block1a104.port_b_data_out_clock = "clock1";
defparam ram_block1a104.port_b_data_width = 1;
defparam ram_block1a104.port_b_first_address = 0;
defparam ram_block1a104.port_b_first_bit_number = 104;
defparam ram_block1a104.port_b_last_address = 7;
defparam ram_block1a104.port_b_logical_ram_depth = 8;
defparam ram_block1a104.port_b_logical_ram_width = 258;
defparam ram_block1a104.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a104.port_b_read_enable_clock = "clock1";
defparam ram_block1a104.ram_block_type = "auto";

cycloneive_ram_block ram_block1a103(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[103]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a103_PORTBDATAOUT_bus));
defparam ram_block1a103.clk1_output_clock_enable = "ena1";
defparam ram_block1a103.data_interleave_offset_in_bits = 1;
defparam ram_block1a103.data_interleave_width_in_bits = 1;
defparam ram_block1a103.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a103.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a103.operation_mode = "dual_port";
defparam ram_block1a103.port_a_address_clear = "none";
defparam ram_block1a103.port_a_address_width = 3;
defparam ram_block1a103.port_a_data_out_clear = "none";
defparam ram_block1a103.port_a_data_out_clock = "none";
defparam ram_block1a103.port_a_data_width = 1;
defparam ram_block1a103.port_a_first_address = 0;
defparam ram_block1a103.port_a_first_bit_number = 103;
defparam ram_block1a103.port_a_last_address = 7;
defparam ram_block1a103.port_a_logical_ram_depth = 8;
defparam ram_block1a103.port_a_logical_ram_width = 258;
defparam ram_block1a103.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a103.port_b_address_clear = "none";
defparam ram_block1a103.port_b_address_clock = "clock1";
defparam ram_block1a103.port_b_address_width = 3;
defparam ram_block1a103.port_b_data_out_clear = "none";
defparam ram_block1a103.port_b_data_out_clock = "clock1";
defparam ram_block1a103.port_b_data_width = 1;
defparam ram_block1a103.port_b_first_address = 0;
defparam ram_block1a103.port_b_first_bit_number = 103;
defparam ram_block1a103.port_b_last_address = 7;
defparam ram_block1a103.port_b_logical_ram_depth = 8;
defparam ram_block1a103.port_b_logical_ram_width = 258;
defparam ram_block1a103.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a103.port_b_read_enable_clock = "clock1";
defparam ram_block1a103.ram_block_type = "auto";

cycloneive_ram_block ram_block1a102(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[102]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a102_PORTBDATAOUT_bus));
defparam ram_block1a102.clk1_output_clock_enable = "ena1";
defparam ram_block1a102.data_interleave_offset_in_bits = 1;
defparam ram_block1a102.data_interleave_width_in_bits = 1;
defparam ram_block1a102.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a102.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a102.operation_mode = "dual_port";
defparam ram_block1a102.port_a_address_clear = "none";
defparam ram_block1a102.port_a_address_width = 3;
defparam ram_block1a102.port_a_data_out_clear = "none";
defparam ram_block1a102.port_a_data_out_clock = "none";
defparam ram_block1a102.port_a_data_width = 1;
defparam ram_block1a102.port_a_first_address = 0;
defparam ram_block1a102.port_a_first_bit_number = 102;
defparam ram_block1a102.port_a_last_address = 7;
defparam ram_block1a102.port_a_logical_ram_depth = 8;
defparam ram_block1a102.port_a_logical_ram_width = 258;
defparam ram_block1a102.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a102.port_b_address_clear = "none";
defparam ram_block1a102.port_b_address_clock = "clock1";
defparam ram_block1a102.port_b_address_width = 3;
defparam ram_block1a102.port_b_data_out_clear = "none";
defparam ram_block1a102.port_b_data_out_clock = "clock1";
defparam ram_block1a102.port_b_data_width = 1;
defparam ram_block1a102.port_b_first_address = 0;
defparam ram_block1a102.port_b_first_bit_number = 102;
defparam ram_block1a102.port_b_last_address = 7;
defparam ram_block1a102.port_b_logical_ram_depth = 8;
defparam ram_block1a102.port_b_logical_ram_width = 258;
defparam ram_block1a102.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a102.port_b_read_enable_clock = "clock1";
defparam ram_block1a102.ram_block_type = "auto";

cycloneive_ram_block ram_block1a101(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[101]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a101_PORTBDATAOUT_bus));
defparam ram_block1a101.clk1_output_clock_enable = "ena1";
defparam ram_block1a101.data_interleave_offset_in_bits = 1;
defparam ram_block1a101.data_interleave_width_in_bits = 1;
defparam ram_block1a101.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a101.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a101.operation_mode = "dual_port";
defparam ram_block1a101.port_a_address_clear = "none";
defparam ram_block1a101.port_a_address_width = 3;
defparam ram_block1a101.port_a_data_out_clear = "none";
defparam ram_block1a101.port_a_data_out_clock = "none";
defparam ram_block1a101.port_a_data_width = 1;
defparam ram_block1a101.port_a_first_address = 0;
defparam ram_block1a101.port_a_first_bit_number = 101;
defparam ram_block1a101.port_a_last_address = 7;
defparam ram_block1a101.port_a_logical_ram_depth = 8;
defparam ram_block1a101.port_a_logical_ram_width = 258;
defparam ram_block1a101.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a101.port_b_address_clear = "none";
defparam ram_block1a101.port_b_address_clock = "clock1";
defparam ram_block1a101.port_b_address_width = 3;
defparam ram_block1a101.port_b_data_out_clear = "none";
defparam ram_block1a101.port_b_data_out_clock = "clock1";
defparam ram_block1a101.port_b_data_width = 1;
defparam ram_block1a101.port_b_first_address = 0;
defparam ram_block1a101.port_b_first_bit_number = 101;
defparam ram_block1a101.port_b_last_address = 7;
defparam ram_block1a101.port_b_logical_ram_depth = 8;
defparam ram_block1a101.port_b_logical_ram_width = 258;
defparam ram_block1a101.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a101.port_b_read_enable_clock = "clock1";
defparam ram_block1a101.ram_block_type = "auto";

cycloneive_ram_block ram_block1a100(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[100]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a100_PORTBDATAOUT_bus));
defparam ram_block1a100.clk1_output_clock_enable = "ena1";
defparam ram_block1a100.data_interleave_offset_in_bits = 1;
defparam ram_block1a100.data_interleave_width_in_bits = 1;
defparam ram_block1a100.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a100.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a100.operation_mode = "dual_port";
defparam ram_block1a100.port_a_address_clear = "none";
defparam ram_block1a100.port_a_address_width = 3;
defparam ram_block1a100.port_a_data_out_clear = "none";
defparam ram_block1a100.port_a_data_out_clock = "none";
defparam ram_block1a100.port_a_data_width = 1;
defparam ram_block1a100.port_a_first_address = 0;
defparam ram_block1a100.port_a_first_bit_number = 100;
defparam ram_block1a100.port_a_last_address = 7;
defparam ram_block1a100.port_a_logical_ram_depth = 8;
defparam ram_block1a100.port_a_logical_ram_width = 258;
defparam ram_block1a100.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a100.port_b_address_clear = "none";
defparam ram_block1a100.port_b_address_clock = "clock1";
defparam ram_block1a100.port_b_address_width = 3;
defparam ram_block1a100.port_b_data_out_clear = "none";
defparam ram_block1a100.port_b_data_out_clock = "clock1";
defparam ram_block1a100.port_b_data_width = 1;
defparam ram_block1a100.port_b_first_address = 0;
defparam ram_block1a100.port_b_first_bit_number = 100;
defparam ram_block1a100.port_b_last_address = 7;
defparam ram_block1a100.port_b_logical_ram_depth = 8;
defparam ram_block1a100.port_b_logical_ram_width = 258;
defparam ram_block1a100.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a100.port_b_read_enable_clock = "clock1";
defparam ram_block1a100.ram_block_type = "auto";

cycloneive_ram_block ram_block1a234(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[234]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a234_PORTBDATAOUT_bus));
defparam ram_block1a234.clk1_output_clock_enable = "ena1";
defparam ram_block1a234.data_interleave_offset_in_bits = 1;
defparam ram_block1a234.data_interleave_width_in_bits = 1;
defparam ram_block1a234.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a234.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a234.operation_mode = "dual_port";
defparam ram_block1a234.port_a_address_clear = "none";
defparam ram_block1a234.port_a_address_width = 3;
defparam ram_block1a234.port_a_data_out_clear = "none";
defparam ram_block1a234.port_a_data_out_clock = "none";
defparam ram_block1a234.port_a_data_width = 1;
defparam ram_block1a234.port_a_first_address = 0;
defparam ram_block1a234.port_a_first_bit_number = 234;
defparam ram_block1a234.port_a_last_address = 7;
defparam ram_block1a234.port_a_logical_ram_depth = 8;
defparam ram_block1a234.port_a_logical_ram_width = 258;
defparam ram_block1a234.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a234.port_b_address_clear = "none";
defparam ram_block1a234.port_b_address_clock = "clock1";
defparam ram_block1a234.port_b_address_width = 3;
defparam ram_block1a234.port_b_data_out_clear = "none";
defparam ram_block1a234.port_b_data_out_clock = "clock1";
defparam ram_block1a234.port_b_data_width = 1;
defparam ram_block1a234.port_b_first_address = 0;
defparam ram_block1a234.port_b_first_bit_number = 234;
defparam ram_block1a234.port_b_last_address = 7;
defparam ram_block1a234.port_b_logical_ram_depth = 8;
defparam ram_block1a234.port_b_logical_ram_width = 258;
defparam ram_block1a234.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a234.port_b_read_enable_clock = "clock1";
defparam ram_block1a234.ram_block_type = "auto";

cycloneive_ram_block ram_block1a233(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[233]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a233_PORTBDATAOUT_bus));
defparam ram_block1a233.clk1_output_clock_enable = "ena1";
defparam ram_block1a233.data_interleave_offset_in_bits = 1;
defparam ram_block1a233.data_interleave_width_in_bits = 1;
defparam ram_block1a233.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a233.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a233.operation_mode = "dual_port";
defparam ram_block1a233.port_a_address_clear = "none";
defparam ram_block1a233.port_a_address_width = 3;
defparam ram_block1a233.port_a_data_out_clear = "none";
defparam ram_block1a233.port_a_data_out_clock = "none";
defparam ram_block1a233.port_a_data_width = 1;
defparam ram_block1a233.port_a_first_address = 0;
defparam ram_block1a233.port_a_first_bit_number = 233;
defparam ram_block1a233.port_a_last_address = 7;
defparam ram_block1a233.port_a_logical_ram_depth = 8;
defparam ram_block1a233.port_a_logical_ram_width = 258;
defparam ram_block1a233.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a233.port_b_address_clear = "none";
defparam ram_block1a233.port_b_address_clock = "clock1";
defparam ram_block1a233.port_b_address_width = 3;
defparam ram_block1a233.port_b_data_out_clear = "none";
defparam ram_block1a233.port_b_data_out_clock = "clock1";
defparam ram_block1a233.port_b_data_width = 1;
defparam ram_block1a233.port_b_first_address = 0;
defparam ram_block1a233.port_b_first_bit_number = 233;
defparam ram_block1a233.port_b_last_address = 7;
defparam ram_block1a233.port_b_logical_ram_depth = 8;
defparam ram_block1a233.port_b_logical_ram_width = 258;
defparam ram_block1a233.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a233.port_b_read_enable_clock = "clock1";
defparam ram_block1a233.ram_block_type = "auto";

cycloneive_ram_block ram_block1a232(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[232]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a232_PORTBDATAOUT_bus));
defparam ram_block1a232.clk1_output_clock_enable = "ena1";
defparam ram_block1a232.data_interleave_offset_in_bits = 1;
defparam ram_block1a232.data_interleave_width_in_bits = 1;
defparam ram_block1a232.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a232.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a232.operation_mode = "dual_port";
defparam ram_block1a232.port_a_address_clear = "none";
defparam ram_block1a232.port_a_address_width = 3;
defparam ram_block1a232.port_a_data_out_clear = "none";
defparam ram_block1a232.port_a_data_out_clock = "none";
defparam ram_block1a232.port_a_data_width = 1;
defparam ram_block1a232.port_a_first_address = 0;
defparam ram_block1a232.port_a_first_bit_number = 232;
defparam ram_block1a232.port_a_last_address = 7;
defparam ram_block1a232.port_a_logical_ram_depth = 8;
defparam ram_block1a232.port_a_logical_ram_width = 258;
defparam ram_block1a232.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a232.port_b_address_clear = "none";
defparam ram_block1a232.port_b_address_clock = "clock1";
defparam ram_block1a232.port_b_address_width = 3;
defparam ram_block1a232.port_b_data_out_clear = "none";
defparam ram_block1a232.port_b_data_out_clock = "clock1";
defparam ram_block1a232.port_b_data_width = 1;
defparam ram_block1a232.port_b_first_address = 0;
defparam ram_block1a232.port_b_first_bit_number = 232;
defparam ram_block1a232.port_b_last_address = 7;
defparam ram_block1a232.port_b_logical_ram_depth = 8;
defparam ram_block1a232.port_b_logical_ram_width = 258;
defparam ram_block1a232.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a232.port_b_read_enable_clock = "clock1";
defparam ram_block1a232.ram_block_type = "auto";

cycloneive_ram_block ram_block1a231(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[231]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a231_PORTBDATAOUT_bus));
defparam ram_block1a231.clk1_output_clock_enable = "ena1";
defparam ram_block1a231.data_interleave_offset_in_bits = 1;
defparam ram_block1a231.data_interleave_width_in_bits = 1;
defparam ram_block1a231.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a231.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a231.operation_mode = "dual_port";
defparam ram_block1a231.port_a_address_clear = "none";
defparam ram_block1a231.port_a_address_width = 3;
defparam ram_block1a231.port_a_data_out_clear = "none";
defparam ram_block1a231.port_a_data_out_clock = "none";
defparam ram_block1a231.port_a_data_width = 1;
defparam ram_block1a231.port_a_first_address = 0;
defparam ram_block1a231.port_a_first_bit_number = 231;
defparam ram_block1a231.port_a_last_address = 7;
defparam ram_block1a231.port_a_logical_ram_depth = 8;
defparam ram_block1a231.port_a_logical_ram_width = 258;
defparam ram_block1a231.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a231.port_b_address_clear = "none";
defparam ram_block1a231.port_b_address_clock = "clock1";
defparam ram_block1a231.port_b_address_width = 3;
defparam ram_block1a231.port_b_data_out_clear = "none";
defparam ram_block1a231.port_b_data_out_clock = "clock1";
defparam ram_block1a231.port_b_data_width = 1;
defparam ram_block1a231.port_b_first_address = 0;
defparam ram_block1a231.port_b_first_bit_number = 231;
defparam ram_block1a231.port_b_last_address = 7;
defparam ram_block1a231.port_b_logical_ram_depth = 8;
defparam ram_block1a231.port_b_logical_ram_width = 258;
defparam ram_block1a231.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a231.port_b_read_enable_clock = "clock1";
defparam ram_block1a231.ram_block_type = "auto";

cycloneive_ram_block ram_block1a230(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[230]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a230_PORTBDATAOUT_bus));
defparam ram_block1a230.clk1_output_clock_enable = "ena1";
defparam ram_block1a230.data_interleave_offset_in_bits = 1;
defparam ram_block1a230.data_interleave_width_in_bits = 1;
defparam ram_block1a230.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a230.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a230.operation_mode = "dual_port";
defparam ram_block1a230.port_a_address_clear = "none";
defparam ram_block1a230.port_a_address_width = 3;
defparam ram_block1a230.port_a_data_out_clear = "none";
defparam ram_block1a230.port_a_data_out_clock = "none";
defparam ram_block1a230.port_a_data_width = 1;
defparam ram_block1a230.port_a_first_address = 0;
defparam ram_block1a230.port_a_first_bit_number = 230;
defparam ram_block1a230.port_a_last_address = 7;
defparam ram_block1a230.port_a_logical_ram_depth = 8;
defparam ram_block1a230.port_a_logical_ram_width = 258;
defparam ram_block1a230.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a230.port_b_address_clear = "none";
defparam ram_block1a230.port_b_address_clock = "clock1";
defparam ram_block1a230.port_b_address_width = 3;
defparam ram_block1a230.port_b_data_out_clear = "none";
defparam ram_block1a230.port_b_data_out_clock = "clock1";
defparam ram_block1a230.port_b_data_width = 1;
defparam ram_block1a230.port_b_first_address = 0;
defparam ram_block1a230.port_b_first_bit_number = 230;
defparam ram_block1a230.port_b_last_address = 7;
defparam ram_block1a230.port_b_logical_ram_depth = 8;
defparam ram_block1a230.port_b_logical_ram_width = 258;
defparam ram_block1a230.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a230.port_b_read_enable_clock = "clock1";
defparam ram_block1a230.ram_block_type = "auto";

cycloneive_ram_block ram_block1a229(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[229]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a229_PORTBDATAOUT_bus));
defparam ram_block1a229.clk1_output_clock_enable = "ena1";
defparam ram_block1a229.data_interleave_offset_in_bits = 1;
defparam ram_block1a229.data_interleave_width_in_bits = 1;
defparam ram_block1a229.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a229.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a229.operation_mode = "dual_port";
defparam ram_block1a229.port_a_address_clear = "none";
defparam ram_block1a229.port_a_address_width = 3;
defparam ram_block1a229.port_a_data_out_clear = "none";
defparam ram_block1a229.port_a_data_out_clock = "none";
defparam ram_block1a229.port_a_data_width = 1;
defparam ram_block1a229.port_a_first_address = 0;
defparam ram_block1a229.port_a_first_bit_number = 229;
defparam ram_block1a229.port_a_last_address = 7;
defparam ram_block1a229.port_a_logical_ram_depth = 8;
defparam ram_block1a229.port_a_logical_ram_width = 258;
defparam ram_block1a229.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a229.port_b_address_clear = "none";
defparam ram_block1a229.port_b_address_clock = "clock1";
defparam ram_block1a229.port_b_address_width = 3;
defparam ram_block1a229.port_b_data_out_clear = "none";
defparam ram_block1a229.port_b_data_out_clock = "clock1";
defparam ram_block1a229.port_b_data_width = 1;
defparam ram_block1a229.port_b_first_address = 0;
defparam ram_block1a229.port_b_first_bit_number = 229;
defparam ram_block1a229.port_b_last_address = 7;
defparam ram_block1a229.port_b_logical_ram_depth = 8;
defparam ram_block1a229.port_b_logical_ram_width = 258;
defparam ram_block1a229.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a229.port_b_read_enable_clock = "clock1";
defparam ram_block1a229.ram_block_type = "auto";

cycloneive_ram_block ram_block1a228(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[228]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a228_PORTBDATAOUT_bus));
defparam ram_block1a228.clk1_output_clock_enable = "ena1";
defparam ram_block1a228.data_interleave_offset_in_bits = 1;
defparam ram_block1a228.data_interleave_width_in_bits = 1;
defparam ram_block1a228.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a228.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a228.operation_mode = "dual_port";
defparam ram_block1a228.port_a_address_clear = "none";
defparam ram_block1a228.port_a_address_width = 3;
defparam ram_block1a228.port_a_data_out_clear = "none";
defparam ram_block1a228.port_a_data_out_clock = "none";
defparam ram_block1a228.port_a_data_width = 1;
defparam ram_block1a228.port_a_first_address = 0;
defparam ram_block1a228.port_a_first_bit_number = 228;
defparam ram_block1a228.port_a_last_address = 7;
defparam ram_block1a228.port_a_logical_ram_depth = 8;
defparam ram_block1a228.port_a_logical_ram_width = 258;
defparam ram_block1a228.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a228.port_b_address_clear = "none";
defparam ram_block1a228.port_b_address_clock = "clock1";
defparam ram_block1a228.port_b_address_width = 3;
defparam ram_block1a228.port_b_data_out_clear = "none";
defparam ram_block1a228.port_b_data_out_clock = "clock1";
defparam ram_block1a228.port_b_data_width = 1;
defparam ram_block1a228.port_b_first_address = 0;
defparam ram_block1a228.port_b_first_bit_number = 228;
defparam ram_block1a228.port_b_last_address = 7;
defparam ram_block1a228.port_b_logical_ram_depth = 8;
defparam ram_block1a228.port_b_logical_ram_width = 258;
defparam ram_block1a228.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a228.port_b_read_enable_clock = "clock1";
defparam ram_block1a228.ram_block_type = "auto";

cycloneive_ram_block ram_block1a42(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[42]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a42_PORTBDATAOUT_bus));
defparam ram_block1a42.clk1_output_clock_enable = "ena1";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a42.operation_mode = "dual_port";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 3;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "none";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 0;
defparam ram_block1a42.port_a_first_bit_number = 42;
defparam ram_block1a42.port_a_last_address = 7;
defparam ram_block1a42.port_a_logical_ram_depth = 8;
defparam ram_block1a42.port_a_logical_ram_width = 258;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a42.port_b_address_clear = "none";
defparam ram_block1a42.port_b_address_clock = "clock1";
defparam ram_block1a42.port_b_address_width = 3;
defparam ram_block1a42.port_b_data_out_clear = "none";
defparam ram_block1a42.port_b_data_out_clock = "clock1";
defparam ram_block1a42.port_b_data_width = 1;
defparam ram_block1a42.port_b_first_address = 0;
defparam ram_block1a42.port_b_first_bit_number = 42;
defparam ram_block1a42.port_b_last_address = 7;
defparam ram_block1a42.port_b_logical_ram_depth = 8;
defparam ram_block1a42.port_b_logical_ram_width = 258;
defparam ram_block1a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a42.port_b_read_enable_clock = "clock1";
defparam ram_block1a42.ram_block_type = "auto";

cycloneive_ram_block ram_block1a41(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[41]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a41_PORTBDATAOUT_bus));
defparam ram_block1a41.clk1_output_clock_enable = "ena1";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a41.operation_mode = "dual_port";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 3;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "none";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 0;
defparam ram_block1a41.port_a_first_bit_number = 41;
defparam ram_block1a41.port_a_last_address = 7;
defparam ram_block1a41.port_a_logical_ram_depth = 8;
defparam ram_block1a41.port_a_logical_ram_width = 258;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a41.port_b_address_clear = "none";
defparam ram_block1a41.port_b_address_clock = "clock1";
defparam ram_block1a41.port_b_address_width = 3;
defparam ram_block1a41.port_b_data_out_clear = "none";
defparam ram_block1a41.port_b_data_out_clock = "clock1";
defparam ram_block1a41.port_b_data_width = 1;
defparam ram_block1a41.port_b_first_address = 0;
defparam ram_block1a41.port_b_first_bit_number = 41;
defparam ram_block1a41.port_b_last_address = 7;
defparam ram_block1a41.port_b_logical_ram_depth = 8;
defparam ram_block1a41.port_b_logical_ram_width = 258;
defparam ram_block1a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a41.port_b_read_enable_clock = "clock1";
defparam ram_block1a41.ram_block_type = "auto";

cycloneive_ram_block ram_block1a40(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[40]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a40_PORTBDATAOUT_bus));
defparam ram_block1a40.clk1_output_clock_enable = "ena1";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a40.operation_mode = "dual_port";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 3;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "none";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 0;
defparam ram_block1a40.port_a_first_bit_number = 40;
defparam ram_block1a40.port_a_last_address = 7;
defparam ram_block1a40.port_a_logical_ram_depth = 8;
defparam ram_block1a40.port_a_logical_ram_width = 258;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a40.port_b_address_clear = "none";
defparam ram_block1a40.port_b_address_clock = "clock1";
defparam ram_block1a40.port_b_address_width = 3;
defparam ram_block1a40.port_b_data_out_clear = "none";
defparam ram_block1a40.port_b_data_out_clock = "clock1";
defparam ram_block1a40.port_b_data_width = 1;
defparam ram_block1a40.port_b_first_address = 0;
defparam ram_block1a40.port_b_first_bit_number = 40;
defparam ram_block1a40.port_b_last_address = 7;
defparam ram_block1a40.port_b_logical_ram_depth = 8;
defparam ram_block1a40.port_b_logical_ram_width = 258;
defparam ram_block1a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a40.port_b_read_enable_clock = "clock1";
defparam ram_block1a40.ram_block_type = "auto";

cycloneive_ram_block ram_block1a39(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[39]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a39_PORTBDATAOUT_bus));
defparam ram_block1a39.clk1_output_clock_enable = "ena1";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a39.operation_mode = "dual_port";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 3;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "none";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 0;
defparam ram_block1a39.port_a_first_bit_number = 39;
defparam ram_block1a39.port_a_last_address = 7;
defparam ram_block1a39.port_a_logical_ram_depth = 8;
defparam ram_block1a39.port_a_logical_ram_width = 258;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a39.port_b_address_clear = "none";
defparam ram_block1a39.port_b_address_clock = "clock1";
defparam ram_block1a39.port_b_address_width = 3;
defparam ram_block1a39.port_b_data_out_clear = "none";
defparam ram_block1a39.port_b_data_out_clock = "clock1";
defparam ram_block1a39.port_b_data_width = 1;
defparam ram_block1a39.port_b_first_address = 0;
defparam ram_block1a39.port_b_first_bit_number = 39;
defparam ram_block1a39.port_b_last_address = 7;
defparam ram_block1a39.port_b_logical_ram_depth = 8;
defparam ram_block1a39.port_b_logical_ram_width = 258;
defparam ram_block1a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a39.port_b_read_enable_clock = "clock1";
defparam ram_block1a39.ram_block_type = "auto";

cycloneive_ram_block ram_block1a38(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[38]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a38_PORTBDATAOUT_bus));
defparam ram_block1a38.clk1_output_clock_enable = "ena1";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a38.operation_mode = "dual_port";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 3;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "none";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 0;
defparam ram_block1a38.port_a_first_bit_number = 38;
defparam ram_block1a38.port_a_last_address = 7;
defparam ram_block1a38.port_a_logical_ram_depth = 8;
defparam ram_block1a38.port_a_logical_ram_width = 258;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a38.port_b_address_clear = "none";
defparam ram_block1a38.port_b_address_clock = "clock1";
defparam ram_block1a38.port_b_address_width = 3;
defparam ram_block1a38.port_b_data_out_clear = "none";
defparam ram_block1a38.port_b_data_out_clock = "clock1";
defparam ram_block1a38.port_b_data_width = 1;
defparam ram_block1a38.port_b_first_address = 0;
defparam ram_block1a38.port_b_first_bit_number = 38;
defparam ram_block1a38.port_b_last_address = 7;
defparam ram_block1a38.port_b_logical_ram_depth = 8;
defparam ram_block1a38.port_b_logical_ram_width = 258;
defparam ram_block1a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a38.port_b_read_enable_clock = "clock1";
defparam ram_block1a38.ram_block_type = "auto";

cycloneive_ram_block ram_block1a37(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[37]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a37_PORTBDATAOUT_bus));
defparam ram_block1a37.clk1_output_clock_enable = "ena1";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a37.operation_mode = "dual_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 3;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 0;
defparam ram_block1a37.port_a_first_bit_number = 37;
defparam ram_block1a37.port_a_last_address = 7;
defparam ram_block1a37.port_a_logical_ram_depth = 8;
defparam ram_block1a37.port_a_logical_ram_width = 258;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a37.port_b_address_clear = "none";
defparam ram_block1a37.port_b_address_clock = "clock1";
defparam ram_block1a37.port_b_address_width = 3;
defparam ram_block1a37.port_b_data_out_clear = "none";
defparam ram_block1a37.port_b_data_out_clock = "clock1";
defparam ram_block1a37.port_b_data_width = 1;
defparam ram_block1a37.port_b_first_address = 0;
defparam ram_block1a37.port_b_first_bit_number = 37;
defparam ram_block1a37.port_b_last_address = 7;
defparam ram_block1a37.port_b_logical_ram_depth = 8;
defparam ram_block1a37.port_b_logical_ram_width = 258;
defparam ram_block1a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a37.port_b_read_enable_clock = "clock1";
defparam ram_block1a37.ram_block_type = "auto";

cycloneive_ram_block ram_block1a36(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[36]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a36_PORTBDATAOUT_bus));
defparam ram_block1a36.clk1_output_clock_enable = "ena1";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a36.operation_mode = "dual_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 3;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 0;
defparam ram_block1a36.port_a_first_bit_number = 36;
defparam ram_block1a36.port_a_last_address = 7;
defparam ram_block1a36.port_a_logical_ram_depth = 8;
defparam ram_block1a36.port_a_logical_ram_width = 258;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a36.port_b_address_clear = "none";
defparam ram_block1a36.port_b_address_clock = "clock1";
defparam ram_block1a36.port_b_address_width = 3;
defparam ram_block1a36.port_b_data_out_clear = "none";
defparam ram_block1a36.port_b_data_out_clock = "clock1";
defparam ram_block1a36.port_b_data_width = 1;
defparam ram_block1a36.port_b_first_address = 0;
defparam ram_block1a36.port_b_first_bit_number = 36;
defparam ram_block1a36.port_b_last_address = 7;
defparam ram_block1a36.port_b_logical_ram_depth = 8;
defparam ram_block1a36.port_b_logical_ram_width = 258;
defparam ram_block1a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a36.port_b_read_enable_clock = "clock1";
defparam ram_block1a36.ram_block_type = "auto";

cycloneive_ram_block ram_block1a186(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[186]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a186_PORTBDATAOUT_bus));
defparam ram_block1a186.clk1_output_clock_enable = "ena1";
defparam ram_block1a186.data_interleave_offset_in_bits = 1;
defparam ram_block1a186.data_interleave_width_in_bits = 1;
defparam ram_block1a186.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a186.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a186.operation_mode = "dual_port";
defparam ram_block1a186.port_a_address_clear = "none";
defparam ram_block1a186.port_a_address_width = 3;
defparam ram_block1a186.port_a_data_out_clear = "none";
defparam ram_block1a186.port_a_data_out_clock = "none";
defparam ram_block1a186.port_a_data_width = 1;
defparam ram_block1a186.port_a_first_address = 0;
defparam ram_block1a186.port_a_first_bit_number = 186;
defparam ram_block1a186.port_a_last_address = 7;
defparam ram_block1a186.port_a_logical_ram_depth = 8;
defparam ram_block1a186.port_a_logical_ram_width = 258;
defparam ram_block1a186.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a186.port_b_address_clear = "none";
defparam ram_block1a186.port_b_address_clock = "clock1";
defparam ram_block1a186.port_b_address_width = 3;
defparam ram_block1a186.port_b_data_out_clear = "none";
defparam ram_block1a186.port_b_data_out_clock = "clock1";
defparam ram_block1a186.port_b_data_width = 1;
defparam ram_block1a186.port_b_first_address = 0;
defparam ram_block1a186.port_b_first_bit_number = 186;
defparam ram_block1a186.port_b_last_address = 7;
defparam ram_block1a186.port_b_logical_ram_depth = 8;
defparam ram_block1a186.port_b_logical_ram_width = 258;
defparam ram_block1a186.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a186.port_b_read_enable_clock = "clock1";
defparam ram_block1a186.ram_block_type = "auto";

cycloneive_ram_block ram_block1a185(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[185]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a185_PORTBDATAOUT_bus));
defparam ram_block1a185.clk1_output_clock_enable = "ena1";
defparam ram_block1a185.data_interleave_offset_in_bits = 1;
defparam ram_block1a185.data_interleave_width_in_bits = 1;
defparam ram_block1a185.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a185.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a185.operation_mode = "dual_port";
defparam ram_block1a185.port_a_address_clear = "none";
defparam ram_block1a185.port_a_address_width = 3;
defparam ram_block1a185.port_a_data_out_clear = "none";
defparam ram_block1a185.port_a_data_out_clock = "none";
defparam ram_block1a185.port_a_data_width = 1;
defparam ram_block1a185.port_a_first_address = 0;
defparam ram_block1a185.port_a_first_bit_number = 185;
defparam ram_block1a185.port_a_last_address = 7;
defparam ram_block1a185.port_a_logical_ram_depth = 8;
defparam ram_block1a185.port_a_logical_ram_width = 258;
defparam ram_block1a185.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a185.port_b_address_clear = "none";
defparam ram_block1a185.port_b_address_clock = "clock1";
defparam ram_block1a185.port_b_address_width = 3;
defparam ram_block1a185.port_b_data_out_clear = "none";
defparam ram_block1a185.port_b_data_out_clock = "clock1";
defparam ram_block1a185.port_b_data_width = 1;
defparam ram_block1a185.port_b_first_address = 0;
defparam ram_block1a185.port_b_first_bit_number = 185;
defparam ram_block1a185.port_b_last_address = 7;
defparam ram_block1a185.port_b_logical_ram_depth = 8;
defparam ram_block1a185.port_b_logical_ram_width = 258;
defparam ram_block1a185.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a185.port_b_read_enable_clock = "clock1";
defparam ram_block1a185.ram_block_type = "auto";

cycloneive_ram_block ram_block1a184(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[184]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a184_PORTBDATAOUT_bus));
defparam ram_block1a184.clk1_output_clock_enable = "ena1";
defparam ram_block1a184.data_interleave_offset_in_bits = 1;
defparam ram_block1a184.data_interleave_width_in_bits = 1;
defparam ram_block1a184.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a184.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a184.operation_mode = "dual_port";
defparam ram_block1a184.port_a_address_clear = "none";
defparam ram_block1a184.port_a_address_width = 3;
defparam ram_block1a184.port_a_data_out_clear = "none";
defparam ram_block1a184.port_a_data_out_clock = "none";
defparam ram_block1a184.port_a_data_width = 1;
defparam ram_block1a184.port_a_first_address = 0;
defparam ram_block1a184.port_a_first_bit_number = 184;
defparam ram_block1a184.port_a_last_address = 7;
defparam ram_block1a184.port_a_logical_ram_depth = 8;
defparam ram_block1a184.port_a_logical_ram_width = 258;
defparam ram_block1a184.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a184.port_b_address_clear = "none";
defparam ram_block1a184.port_b_address_clock = "clock1";
defparam ram_block1a184.port_b_address_width = 3;
defparam ram_block1a184.port_b_data_out_clear = "none";
defparam ram_block1a184.port_b_data_out_clock = "clock1";
defparam ram_block1a184.port_b_data_width = 1;
defparam ram_block1a184.port_b_first_address = 0;
defparam ram_block1a184.port_b_first_bit_number = 184;
defparam ram_block1a184.port_b_last_address = 7;
defparam ram_block1a184.port_b_logical_ram_depth = 8;
defparam ram_block1a184.port_b_logical_ram_width = 258;
defparam ram_block1a184.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a184.port_b_read_enable_clock = "clock1";
defparam ram_block1a184.ram_block_type = "auto";

cycloneive_ram_block ram_block1a183(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[183]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a183_PORTBDATAOUT_bus));
defparam ram_block1a183.clk1_output_clock_enable = "ena1";
defparam ram_block1a183.data_interleave_offset_in_bits = 1;
defparam ram_block1a183.data_interleave_width_in_bits = 1;
defparam ram_block1a183.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a183.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a183.operation_mode = "dual_port";
defparam ram_block1a183.port_a_address_clear = "none";
defparam ram_block1a183.port_a_address_width = 3;
defparam ram_block1a183.port_a_data_out_clear = "none";
defparam ram_block1a183.port_a_data_out_clock = "none";
defparam ram_block1a183.port_a_data_width = 1;
defparam ram_block1a183.port_a_first_address = 0;
defparam ram_block1a183.port_a_first_bit_number = 183;
defparam ram_block1a183.port_a_last_address = 7;
defparam ram_block1a183.port_a_logical_ram_depth = 8;
defparam ram_block1a183.port_a_logical_ram_width = 258;
defparam ram_block1a183.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a183.port_b_address_clear = "none";
defparam ram_block1a183.port_b_address_clock = "clock1";
defparam ram_block1a183.port_b_address_width = 3;
defparam ram_block1a183.port_b_data_out_clear = "none";
defparam ram_block1a183.port_b_data_out_clock = "clock1";
defparam ram_block1a183.port_b_data_width = 1;
defparam ram_block1a183.port_b_first_address = 0;
defparam ram_block1a183.port_b_first_bit_number = 183;
defparam ram_block1a183.port_b_last_address = 7;
defparam ram_block1a183.port_b_logical_ram_depth = 8;
defparam ram_block1a183.port_b_logical_ram_width = 258;
defparam ram_block1a183.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a183.port_b_read_enable_clock = "clock1";
defparam ram_block1a183.ram_block_type = "auto";

cycloneive_ram_block ram_block1a182(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[182]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a182_PORTBDATAOUT_bus));
defparam ram_block1a182.clk1_output_clock_enable = "ena1";
defparam ram_block1a182.data_interleave_offset_in_bits = 1;
defparam ram_block1a182.data_interleave_width_in_bits = 1;
defparam ram_block1a182.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a182.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a182.operation_mode = "dual_port";
defparam ram_block1a182.port_a_address_clear = "none";
defparam ram_block1a182.port_a_address_width = 3;
defparam ram_block1a182.port_a_data_out_clear = "none";
defparam ram_block1a182.port_a_data_out_clock = "none";
defparam ram_block1a182.port_a_data_width = 1;
defparam ram_block1a182.port_a_first_address = 0;
defparam ram_block1a182.port_a_first_bit_number = 182;
defparam ram_block1a182.port_a_last_address = 7;
defparam ram_block1a182.port_a_logical_ram_depth = 8;
defparam ram_block1a182.port_a_logical_ram_width = 258;
defparam ram_block1a182.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a182.port_b_address_clear = "none";
defparam ram_block1a182.port_b_address_clock = "clock1";
defparam ram_block1a182.port_b_address_width = 3;
defparam ram_block1a182.port_b_data_out_clear = "none";
defparam ram_block1a182.port_b_data_out_clock = "clock1";
defparam ram_block1a182.port_b_data_width = 1;
defparam ram_block1a182.port_b_first_address = 0;
defparam ram_block1a182.port_b_first_bit_number = 182;
defparam ram_block1a182.port_b_last_address = 7;
defparam ram_block1a182.port_b_logical_ram_depth = 8;
defparam ram_block1a182.port_b_logical_ram_width = 258;
defparam ram_block1a182.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a182.port_b_read_enable_clock = "clock1";
defparam ram_block1a182.ram_block_type = "auto";

cycloneive_ram_block ram_block1a181(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[181]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a181_PORTBDATAOUT_bus));
defparam ram_block1a181.clk1_output_clock_enable = "ena1";
defparam ram_block1a181.data_interleave_offset_in_bits = 1;
defparam ram_block1a181.data_interleave_width_in_bits = 1;
defparam ram_block1a181.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a181.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a181.operation_mode = "dual_port";
defparam ram_block1a181.port_a_address_clear = "none";
defparam ram_block1a181.port_a_address_width = 3;
defparam ram_block1a181.port_a_data_out_clear = "none";
defparam ram_block1a181.port_a_data_out_clock = "none";
defparam ram_block1a181.port_a_data_width = 1;
defparam ram_block1a181.port_a_first_address = 0;
defparam ram_block1a181.port_a_first_bit_number = 181;
defparam ram_block1a181.port_a_last_address = 7;
defparam ram_block1a181.port_a_logical_ram_depth = 8;
defparam ram_block1a181.port_a_logical_ram_width = 258;
defparam ram_block1a181.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a181.port_b_address_clear = "none";
defparam ram_block1a181.port_b_address_clock = "clock1";
defparam ram_block1a181.port_b_address_width = 3;
defparam ram_block1a181.port_b_data_out_clear = "none";
defparam ram_block1a181.port_b_data_out_clock = "clock1";
defparam ram_block1a181.port_b_data_width = 1;
defparam ram_block1a181.port_b_first_address = 0;
defparam ram_block1a181.port_b_first_bit_number = 181;
defparam ram_block1a181.port_b_last_address = 7;
defparam ram_block1a181.port_b_logical_ram_depth = 8;
defparam ram_block1a181.port_b_logical_ram_width = 258;
defparam ram_block1a181.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a181.port_b_read_enable_clock = "clock1";
defparam ram_block1a181.ram_block_type = "auto";

cycloneive_ram_block ram_block1a180(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[180]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a180_PORTBDATAOUT_bus));
defparam ram_block1a180.clk1_output_clock_enable = "ena1";
defparam ram_block1a180.data_interleave_offset_in_bits = 1;
defparam ram_block1a180.data_interleave_width_in_bits = 1;
defparam ram_block1a180.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a180.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a180.operation_mode = "dual_port";
defparam ram_block1a180.port_a_address_clear = "none";
defparam ram_block1a180.port_a_address_width = 3;
defparam ram_block1a180.port_a_data_out_clear = "none";
defparam ram_block1a180.port_a_data_out_clock = "none";
defparam ram_block1a180.port_a_data_width = 1;
defparam ram_block1a180.port_a_first_address = 0;
defparam ram_block1a180.port_a_first_bit_number = 180;
defparam ram_block1a180.port_a_last_address = 7;
defparam ram_block1a180.port_a_logical_ram_depth = 8;
defparam ram_block1a180.port_a_logical_ram_width = 258;
defparam ram_block1a180.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a180.port_b_address_clear = "none";
defparam ram_block1a180.port_b_address_clock = "clock1";
defparam ram_block1a180.port_b_address_width = 3;
defparam ram_block1a180.port_b_data_out_clear = "none";
defparam ram_block1a180.port_b_data_out_clock = "clock1";
defparam ram_block1a180.port_b_data_width = 1;
defparam ram_block1a180.port_b_first_address = 0;
defparam ram_block1a180.port_b_first_bit_number = 180;
defparam ram_block1a180.port_b_last_address = 7;
defparam ram_block1a180.port_b_logical_ram_depth = 8;
defparam ram_block1a180.port_b_logical_ram_width = 258;
defparam ram_block1a180.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a180.port_b_read_enable_clock = "clock1";
defparam ram_block1a180.ram_block_type = "auto";

cycloneive_ram_block ram_block1a122(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[122]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a122_PORTBDATAOUT_bus));
defparam ram_block1a122.clk1_output_clock_enable = "ena1";
defparam ram_block1a122.data_interleave_offset_in_bits = 1;
defparam ram_block1a122.data_interleave_width_in_bits = 1;
defparam ram_block1a122.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a122.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a122.operation_mode = "dual_port";
defparam ram_block1a122.port_a_address_clear = "none";
defparam ram_block1a122.port_a_address_width = 3;
defparam ram_block1a122.port_a_data_out_clear = "none";
defparam ram_block1a122.port_a_data_out_clock = "none";
defparam ram_block1a122.port_a_data_width = 1;
defparam ram_block1a122.port_a_first_address = 0;
defparam ram_block1a122.port_a_first_bit_number = 122;
defparam ram_block1a122.port_a_last_address = 7;
defparam ram_block1a122.port_a_logical_ram_depth = 8;
defparam ram_block1a122.port_a_logical_ram_width = 258;
defparam ram_block1a122.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a122.port_b_address_clear = "none";
defparam ram_block1a122.port_b_address_clock = "clock1";
defparam ram_block1a122.port_b_address_width = 3;
defparam ram_block1a122.port_b_data_out_clear = "none";
defparam ram_block1a122.port_b_data_out_clock = "clock1";
defparam ram_block1a122.port_b_data_width = 1;
defparam ram_block1a122.port_b_first_address = 0;
defparam ram_block1a122.port_b_first_bit_number = 122;
defparam ram_block1a122.port_b_last_address = 7;
defparam ram_block1a122.port_b_logical_ram_depth = 8;
defparam ram_block1a122.port_b_logical_ram_width = 258;
defparam ram_block1a122.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a122.port_b_read_enable_clock = "clock1";
defparam ram_block1a122.ram_block_type = "auto";

cycloneive_ram_block ram_block1a121(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[121]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a121_PORTBDATAOUT_bus));
defparam ram_block1a121.clk1_output_clock_enable = "ena1";
defparam ram_block1a121.data_interleave_offset_in_bits = 1;
defparam ram_block1a121.data_interleave_width_in_bits = 1;
defparam ram_block1a121.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a121.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a121.operation_mode = "dual_port";
defparam ram_block1a121.port_a_address_clear = "none";
defparam ram_block1a121.port_a_address_width = 3;
defparam ram_block1a121.port_a_data_out_clear = "none";
defparam ram_block1a121.port_a_data_out_clock = "none";
defparam ram_block1a121.port_a_data_width = 1;
defparam ram_block1a121.port_a_first_address = 0;
defparam ram_block1a121.port_a_first_bit_number = 121;
defparam ram_block1a121.port_a_last_address = 7;
defparam ram_block1a121.port_a_logical_ram_depth = 8;
defparam ram_block1a121.port_a_logical_ram_width = 258;
defparam ram_block1a121.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a121.port_b_address_clear = "none";
defparam ram_block1a121.port_b_address_clock = "clock1";
defparam ram_block1a121.port_b_address_width = 3;
defparam ram_block1a121.port_b_data_out_clear = "none";
defparam ram_block1a121.port_b_data_out_clock = "clock1";
defparam ram_block1a121.port_b_data_width = 1;
defparam ram_block1a121.port_b_first_address = 0;
defparam ram_block1a121.port_b_first_bit_number = 121;
defparam ram_block1a121.port_b_last_address = 7;
defparam ram_block1a121.port_b_logical_ram_depth = 8;
defparam ram_block1a121.port_b_logical_ram_width = 258;
defparam ram_block1a121.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a121.port_b_read_enable_clock = "clock1";
defparam ram_block1a121.ram_block_type = "auto";

cycloneive_ram_block ram_block1a120(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[120]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a120_PORTBDATAOUT_bus));
defparam ram_block1a120.clk1_output_clock_enable = "ena1";
defparam ram_block1a120.data_interleave_offset_in_bits = 1;
defparam ram_block1a120.data_interleave_width_in_bits = 1;
defparam ram_block1a120.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a120.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a120.operation_mode = "dual_port";
defparam ram_block1a120.port_a_address_clear = "none";
defparam ram_block1a120.port_a_address_width = 3;
defparam ram_block1a120.port_a_data_out_clear = "none";
defparam ram_block1a120.port_a_data_out_clock = "none";
defparam ram_block1a120.port_a_data_width = 1;
defparam ram_block1a120.port_a_first_address = 0;
defparam ram_block1a120.port_a_first_bit_number = 120;
defparam ram_block1a120.port_a_last_address = 7;
defparam ram_block1a120.port_a_logical_ram_depth = 8;
defparam ram_block1a120.port_a_logical_ram_width = 258;
defparam ram_block1a120.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a120.port_b_address_clear = "none";
defparam ram_block1a120.port_b_address_clock = "clock1";
defparam ram_block1a120.port_b_address_width = 3;
defparam ram_block1a120.port_b_data_out_clear = "none";
defparam ram_block1a120.port_b_data_out_clock = "clock1";
defparam ram_block1a120.port_b_data_width = 1;
defparam ram_block1a120.port_b_first_address = 0;
defparam ram_block1a120.port_b_first_bit_number = 120;
defparam ram_block1a120.port_b_last_address = 7;
defparam ram_block1a120.port_b_logical_ram_depth = 8;
defparam ram_block1a120.port_b_logical_ram_width = 258;
defparam ram_block1a120.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a120.port_b_read_enable_clock = "clock1";
defparam ram_block1a120.ram_block_type = "auto";

cycloneive_ram_block ram_block1a119(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[119]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a119_PORTBDATAOUT_bus));
defparam ram_block1a119.clk1_output_clock_enable = "ena1";
defparam ram_block1a119.data_interleave_offset_in_bits = 1;
defparam ram_block1a119.data_interleave_width_in_bits = 1;
defparam ram_block1a119.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a119.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a119.operation_mode = "dual_port";
defparam ram_block1a119.port_a_address_clear = "none";
defparam ram_block1a119.port_a_address_width = 3;
defparam ram_block1a119.port_a_data_out_clear = "none";
defparam ram_block1a119.port_a_data_out_clock = "none";
defparam ram_block1a119.port_a_data_width = 1;
defparam ram_block1a119.port_a_first_address = 0;
defparam ram_block1a119.port_a_first_bit_number = 119;
defparam ram_block1a119.port_a_last_address = 7;
defparam ram_block1a119.port_a_logical_ram_depth = 8;
defparam ram_block1a119.port_a_logical_ram_width = 258;
defparam ram_block1a119.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a119.port_b_address_clear = "none";
defparam ram_block1a119.port_b_address_clock = "clock1";
defparam ram_block1a119.port_b_address_width = 3;
defparam ram_block1a119.port_b_data_out_clear = "none";
defparam ram_block1a119.port_b_data_out_clock = "clock1";
defparam ram_block1a119.port_b_data_width = 1;
defparam ram_block1a119.port_b_first_address = 0;
defparam ram_block1a119.port_b_first_bit_number = 119;
defparam ram_block1a119.port_b_last_address = 7;
defparam ram_block1a119.port_b_logical_ram_depth = 8;
defparam ram_block1a119.port_b_logical_ram_width = 258;
defparam ram_block1a119.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a119.port_b_read_enable_clock = "clock1";
defparam ram_block1a119.ram_block_type = "auto";

cycloneive_ram_block ram_block1a118(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[118]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a118_PORTBDATAOUT_bus));
defparam ram_block1a118.clk1_output_clock_enable = "ena1";
defparam ram_block1a118.data_interleave_offset_in_bits = 1;
defparam ram_block1a118.data_interleave_width_in_bits = 1;
defparam ram_block1a118.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a118.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a118.operation_mode = "dual_port";
defparam ram_block1a118.port_a_address_clear = "none";
defparam ram_block1a118.port_a_address_width = 3;
defparam ram_block1a118.port_a_data_out_clear = "none";
defparam ram_block1a118.port_a_data_out_clock = "none";
defparam ram_block1a118.port_a_data_width = 1;
defparam ram_block1a118.port_a_first_address = 0;
defparam ram_block1a118.port_a_first_bit_number = 118;
defparam ram_block1a118.port_a_last_address = 7;
defparam ram_block1a118.port_a_logical_ram_depth = 8;
defparam ram_block1a118.port_a_logical_ram_width = 258;
defparam ram_block1a118.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a118.port_b_address_clear = "none";
defparam ram_block1a118.port_b_address_clock = "clock1";
defparam ram_block1a118.port_b_address_width = 3;
defparam ram_block1a118.port_b_data_out_clear = "none";
defparam ram_block1a118.port_b_data_out_clock = "clock1";
defparam ram_block1a118.port_b_data_width = 1;
defparam ram_block1a118.port_b_first_address = 0;
defparam ram_block1a118.port_b_first_bit_number = 118;
defparam ram_block1a118.port_b_last_address = 7;
defparam ram_block1a118.port_b_logical_ram_depth = 8;
defparam ram_block1a118.port_b_logical_ram_width = 258;
defparam ram_block1a118.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a118.port_b_read_enable_clock = "clock1";
defparam ram_block1a118.ram_block_type = "auto";

cycloneive_ram_block ram_block1a117(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[117]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a117_PORTBDATAOUT_bus));
defparam ram_block1a117.clk1_output_clock_enable = "ena1";
defparam ram_block1a117.data_interleave_offset_in_bits = 1;
defparam ram_block1a117.data_interleave_width_in_bits = 1;
defparam ram_block1a117.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a117.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a117.operation_mode = "dual_port";
defparam ram_block1a117.port_a_address_clear = "none";
defparam ram_block1a117.port_a_address_width = 3;
defparam ram_block1a117.port_a_data_out_clear = "none";
defparam ram_block1a117.port_a_data_out_clock = "none";
defparam ram_block1a117.port_a_data_width = 1;
defparam ram_block1a117.port_a_first_address = 0;
defparam ram_block1a117.port_a_first_bit_number = 117;
defparam ram_block1a117.port_a_last_address = 7;
defparam ram_block1a117.port_a_logical_ram_depth = 8;
defparam ram_block1a117.port_a_logical_ram_width = 258;
defparam ram_block1a117.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a117.port_b_address_clear = "none";
defparam ram_block1a117.port_b_address_clock = "clock1";
defparam ram_block1a117.port_b_address_width = 3;
defparam ram_block1a117.port_b_data_out_clear = "none";
defparam ram_block1a117.port_b_data_out_clock = "clock1";
defparam ram_block1a117.port_b_data_width = 1;
defparam ram_block1a117.port_b_first_address = 0;
defparam ram_block1a117.port_b_first_bit_number = 117;
defparam ram_block1a117.port_b_last_address = 7;
defparam ram_block1a117.port_b_logical_ram_depth = 8;
defparam ram_block1a117.port_b_logical_ram_width = 258;
defparam ram_block1a117.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a117.port_b_read_enable_clock = "clock1";
defparam ram_block1a117.ram_block_type = "auto";

cycloneive_ram_block ram_block1a116(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[116]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a116_PORTBDATAOUT_bus));
defparam ram_block1a116.clk1_output_clock_enable = "ena1";
defparam ram_block1a116.data_interleave_offset_in_bits = 1;
defparam ram_block1a116.data_interleave_width_in_bits = 1;
defparam ram_block1a116.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a116.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a116.operation_mode = "dual_port";
defparam ram_block1a116.port_a_address_clear = "none";
defparam ram_block1a116.port_a_address_width = 3;
defparam ram_block1a116.port_a_data_out_clear = "none";
defparam ram_block1a116.port_a_data_out_clock = "none";
defparam ram_block1a116.port_a_data_width = 1;
defparam ram_block1a116.port_a_first_address = 0;
defparam ram_block1a116.port_a_first_bit_number = 116;
defparam ram_block1a116.port_a_last_address = 7;
defparam ram_block1a116.port_a_logical_ram_depth = 8;
defparam ram_block1a116.port_a_logical_ram_width = 258;
defparam ram_block1a116.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a116.port_b_address_clear = "none";
defparam ram_block1a116.port_b_address_clock = "clock1";
defparam ram_block1a116.port_b_address_width = 3;
defparam ram_block1a116.port_b_data_out_clear = "none";
defparam ram_block1a116.port_b_data_out_clock = "clock1";
defparam ram_block1a116.port_b_data_width = 1;
defparam ram_block1a116.port_b_first_address = 0;
defparam ram_block1a116.port_b_first_bit_number = 116;
defparam ram_block1a116.port_b_last_address = 7;
defparam ram_block1a116.port_b_logical_ram_depth = 8;
defparam ram_block1a116.port_b_logical_ram_width = 258;
defparam ram_block1a116.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a116.port_b_read_enable_clock = "clock1";
defparam ram_block1a116.ram_block_type = "auto";

cycloneive_ram_block ram_block1a250(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[250]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a250_PORTBDATAOUT_bus));
defparam ram_block1a250.clk1_output_clock_enable = "ena1";
defparam ram_block1a250.data_interleave_offset_in_bits = 1;
defparam ram_block1a250.data_interleave_width_in_bits = 1;
defparam ram_block1a250.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a250.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a250.operation_mode = "dual_port";
defparam ram_block1a250.port_a_address_clear = "none";
defparam ram_block1a250.port_a_address_width = 3;
defparam ram_block1a250.port_a_data_out_clear = "none";
defparam ram_block1a250.port_a_data_out_clock = "none";
defparam ram_block1a250.port_a_data_width = 1;
defparam ram_block1a250.port_a_first_address = 0;
defparam ram_block1a250.port_a_first_bit_number = 250;
defparam ram_block1a250.port_a_last_address = 7;
defparam ram_block1a250.port_a_logical_ram_depth = 8;
defparam ram_block1a250.port_a_logical_ram_width = 258;
defparam ram_block1a250.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a250.port_b_address_clear = "none";
defparam ram_block1a250.port_b_address_clock = "clock1";
defparam ram_block1a250.port_b_address_width = 3;
defparam ram_block1a250.port_b_data_out_clear = "none";
defparam ram_block1a250.port_b_data_out_clock = "clock1";
defparam ram_block1a250.port_b_data_width = 1;
defparam ram_block1a250.port_b_first_address = 0;
defparam ram_block1a250.port_b_first_bit_number = 250;
defparam ram_block1a250.port_b_last_address = 7;
defparam ram_block1a250.port_b_logical_ram_depth = 8;
defparam ram_block1a250.port_b_logical_ram_width = 258;
defparam ram_block1a250.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a250.port_b_read_enable_clock = "clock1";
defparam ram_block1a250.ram_block_type = "auto";

cycloneive_ram_block ram_block1a249(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[249]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a249_PORTBDATAOUT_bus));
defparam ram_block1a249.clk1_output_clock_enable = "ena1";
defparam ram_block1a249.data_interleave_offset_in_bits = 1;
defparam ram_block1a249.data_interleave_width_in_bits = 1;
defparam ram_block1a249.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a249.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a249.operation_mode = "dual_port";
defparam ram_block1a249.port_a_address_clear = "none";
defparam ram_block1a249.port_a_address_width = 3;
defparam ram_block1a249.port_a_data_out_clear = "none";
defparam ram_block1a249.port_a_data_out_clock = "none";
defparam ram_block1a249.port_a_data_width = 1;
defparam ram_block1a249.port_a_first_address = 0;
defparam ram_block1a249.port_a_first_bit_number = 249;
defparam ram_block1a249.port_a_last_address = 7;
defparam ram_block1a249.port_a_logical_ram_depth = 8;
defparam ram_block1a249.port_a_logical_ram_width = 258;
defparam ram_block1a249.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a249.port_b_address_clear = "none";
defparam ram_block1a249.port_b_address_clock = "clock1";
defparam ram_block1a249.port_b_address_width = 3;
defparam ram_block1a249.port_b_data_out_clear = "none";
defparam ram_block1a249.port_b_data_out_clock = "clock1";
defparam ram_block1a249.port_b_data_width = 1;
defparam ram_block1a249.port_b_first_address = 0;
defparam ram_block1a249.port_b_first_bit_number = 249;
defparam ram_block1a249.port_b_last_address = 7;
defparam ram_block1a249.port_b_logical_ram_depth = 8;
defparam ram_block1a249.port_b_logical_ram_width = 258;
defparam ram_block1a249.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a249.port_b_read_enable_clock = "clock1";
defparam ram_block1a249.ram_block_type = "auto";

cycloneive_ram_block ram_block1a248(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[248]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a248_PORTBDATAOUT_bus));
defparam ram_block1a248.clk1_output_clock_enable = "ena1";
defparam ram_block1a248.data_interleave_offset_in_bits = 1;
defparam ram_block1a248.data_interleave_width_in_bits = 1;
defparam ram_block1a248.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a248.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a248.operation_mode = "dual_port";
defparam ram_block1a248.port_a_address_clear = "none";
defparam ram_block1a248.port_a_address_width = 3;
defparam ram_block1a248.port_a_data_out_clear = "none";
defparam ram_block1a248.port_a_data_out_clock = "none";
defparam ram_block1a248.port_a_data_width = 1;
defparam ram_block1a248.port_a_first_address = 0;
defparam ram_block1a248.port_a_first_bit_number = 248;
defparam ram_block1a248.port_a_last_address = 7;
defparam ram_block1a248.port_a_logical_ram_depth = 8;
defparam ram_block1a248.port_a_logical_ram_width = 258;
defparam ram_block1a248.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a248.port_b_address_clear = "none";
defparam ram_block1a248.port_b_address_clock = "clock1";
defparam ram_block1a248.port_b_address_width = 3;
defparam ram_block1a248.port_b_data_out_clear = "none";
defparam ram_block1a248.port_b_data_out_clock = "clock1";
defparam ram_block1a248.port_b_data_width = 1;
defparam ram_block1a248.port_b_first_address = 0;
defparam ram_block1a248.port_b_first_bit_number = 248;
defparam ram_block1a248.port_b_last_address = 7;
defparam ram_block1a248.port_b_logical_ram_depth = 8;
defparam ram_block1a248.port_b_logical_ram_width = 258;
defparam ram_block1a248.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a248.port_b_read_enable_clock = "clock1";
defparam ram_block1a248.ram_block_type = "auto";

cycloneive_ram_block ram_block1a247(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[247]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a247_PORTBDATAOUT_bus));
defparam ram_block1a247.clk1_output_clock_enable = "ena1";
defparam ram_block1a247.data_interleave_offset_in_bits = 1;
defparam ram_block1a247.data_interleave_width_in_bits = 1;
defparam ram_block1a247.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a247.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a247.operation_mode = "dual_port";
defparam ram_block1a247.port_a_address_clear = "none";
defparam ram_block1a247.port_a_address_width = 3;
defparam ram_block1a247.port_a_data_out_clear = "none";
defparam ram_block1a247.port_a_data_out_clock = "none";
defparam ram_block1a247.port_a_data_width = 1;
defparam ram_block1a247.port_a_first_address = 0;
defparam ram_block1a247.port_a_first_bit_number = 247;
defparam ram_block1a247.port_a_last_address = 7;
defparam ram_block1a247.port_a_logical_ram_depth = 8;
defparam ram_block1a247.port_a_logical_ram_width = 258;
defparam ram_block1a247.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a247.port_b_address_clear = "none";
defparam ram_block1a247.port_b_address_clock = "clock1";
defparam ram_block1a247.port_b_address_width = 3;
defparam ram_block1a247.port_b_data_out_clear = "none";
defparam ram_block1a247.port_b_data_out_clock = "clock1";
defparam ram_block1a247.port_b_data_width = 1;
defparam ram_block1a247.port_b_first_address = 0;
defparam ram_block1a247.port_b_first_bit_number = 247;
defparam ram_block1a247.port_b_last_address = 7;
defparam ram_block1a247.port_b_logical_ram_depth = 8;
defparam ram_block1a247.port_b_logical_ram_width = 258;
defparam ram_block1a247.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a247.port_b_read_enable_clock = "clock1";
defparam ram_block1a247.ram_block_type = "auto";

cycloneive_ram_block ram_block1a246(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[246]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a246_PORTBDATAOUT_bus));
defparam ram_block1a246.clk1_output_clock_enable = "ena1";
defparam ram_block1a246.data_interleave_offset_in_bits = 1;
defparam ram_block1a246.data_interleave_width_in_bits = 1;
defparam ram_block1a246.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a246.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a246.operation_mode = "dual_port";
defparam ram_block1a246.port_a_address_clear = "none";
defparam ram_block1a246.port_a_address_width = 3;
defparam ram_block1a246.port_a_data_out_clear = "none";
defparam ram_block1a246.port_a_data_out_clock = "none";
defparam ram_block1a246.port_a_data_width = 1;
defparam ram_block1a246.port_a_first_address = 0;
defparam ram_block1a246.port_a_first_bit_number = 246;
defparam ram_block1a246.port_a_last_address = 7;
defparam ram_block1a246.port_a_logical_ram_depth = 8;
defparam ram_block1a246.port_a_logical_ram_width = 258;
defparam ram_block1a246.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a246.port_b_address_clear = "none";
defparam ram_block1a246.port_b_address_clock = "clock1";
defparam ram_block1a246.port_b_address_width = 3;
defparam ram_block1a246.port_b_data_out_clear = "none";
defparam ram_block1a246.port_b_data_out_clock = "clock1";
defparam ram_block1a246.port_b_data_width = 1;
defparam ram_block1a246.port_b_first_address = 0;
defparam ram_block1a246.port_b_first_bit_number = 246;
defparam ram_block1a246.port_b_last_address = 7;
defparam ram_block1a246.port_b_logical_ram_depth = 8;
defparam ram_block1a246.port_b_logical_ram_width = 258;
defparam ram_block1a246.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a246.port_b_read_enable_clock = "clock1";
defparam ram_block1a246.ram_block_type = "auto";

cycloneive_ram_block ram_block1a245(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[245]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a245_PORTBDATAOUT_bus));
defparam ram_block1a245.clk1_output_clock_enable = "ena1";
defparam ram_block1a245.data_interleave_offset_in_bits = 1;
defparam ram_block1a245.data_interleave_width_in_bits = 1;
defparam ram_block1a245.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a245.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a245.operation_mode = "dual_port";
defparam ram_block1a245.port_a_address_clear = "none";
defparam ram_block1a245.port_a_address_width = 3;
defparam ram_block1a245.port_a_data_out_clear = "none";
defparam ram_block1a245.port_a_data_out_clock = "none";
defparam ram_block1a245.port_a_data_width = 1;
defparam ram_block1a245.port_a_first_address = 0;
defparam ram_block1a245.port_a_first_bit_number = 245;
defparam ram_block1a245.port_a_last_address = 7;
defparam ram_block1a245.port_a_logical_ram_depth = 8;
defparam ram_block1a245.port_a_logical_ram_width = 258;
defparam ram_block1a245.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a245.port_b_address_clear = "none";
defparam ram_block1a245.port_b_address_clock = "clock1";
defparam ram_block1a245.port_b_address_width = 3;
defparam ram_block1a245.port_b_data_out_clear = "none";
defparam ram_block1a245.port_b_data_out_clock = "clock1";
defparam ram_block1a245.port_b_data_width = 1;
defparam ram_block1a245.port_b_first_address = 0;
defparam ram_block1a245.port_b_first_bit_number = 245;
defparam ram_block1a245.port_b_last_address = 7;
defparam ram_block1a245.port_b_logical_ram_depth = 8;
defparam ram_block1a245.port_b_logical_ram_width = 258;
defparam ram_block1a245.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a245.port_b_read_enable_clock = "clock1";
defparam ram_block1a245.ram_block_type = "auto";

cycloneive_ram_block ram_block1a244(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[244]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a244_PORTBDATAOUT_bus));
defparam ram_block1a244.clk1_output_clock_enable = "ena1";
defparam ram_block1a244.data_interleave_offset_in_bits = 1;
defparam ram_block1a244.data_interleave_width_in_bits = 1;
defparam ram_block1a244.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a244.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a244.operation_mode = "dual_port";
defparam ram_block1a244.port_a_address_clear = "none";
defparam ram_block1a244.port_a_address_width = 3;
defparam ram_block1a244.port_a_data_out_clear = "none";
defparam ram_block1a244.port_a_data_out_clock = "none";
defparam ram_block1a244.port_a_data_width = 1;
defparam ram_block1a244.port_a_first_address = 0;
defparam ram_block1a244.port_a_first_bit_number = 244;
defparam ram_block1a244.port_a_last_address = 7;
defparam ram_block1a244.port_a_logical_ram_depth = 8;
defparam ram_block1a244.port_a_logical_ram_width = 258;
defparam ram_block1a244.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a244.port_b_address_clear = "none";
defparam ram_block1a244.port_b_address_clock = "clock1";
defparam ram_block1a244.port_b_address_width = 3;
defparam ram_block1a244.port_b_data_out_clear = "none";
defparam ram_block1a244.port_b_data_out_clock = "clock1";
defparam ram_block1a244.port_b_data_width = 1;
defparam ram_block1a244.port_b_first_address = 0;
defparam ram_block1a244.port_b_first_bit_number = 244;
defparam ram_block1a244.port_b_last_address = 7;
defparam ram_block1a244.port_b_logical_ram_depth = 8;
defparam ram_block1a244.port_b_logical_ram_width = 258;
defparam ram_block1a244.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a244.port_b_read_enable_clock = "clock1";
defparam ram_block1a244.ram_block_type = "auto";

cycloneive_ram_block ram_block1a58(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[58]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a58_PORTBDATAOUT_bus));
defparam ram_block1a58.clk1_output_clock_enable = "ena1";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a58.operation_mode = "dual_port";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 3;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "none";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 0;
defparam ram_block1a58.port_a_first_bit_number = 58;
defparam ram_block1a58.port_a_last_address = 7;
defparam ram_block1a58.port_a_logical_ram_depth = 8;
defparam ram_block1a58.port_a_logical_ram_width = 258;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a58.port_b_address_clear = "none";
defparam ram_block1a58.port_b_address_clock = "clock1";
defparam ram_block1a58.port_b_address_width = 3;
defparam ram_block1a58.port_b_data_out_clear = "none";
defparam ram_block1a58.port_b_data_out_clock = "clock1";
defparam ram_block1a58.port_b_data_width = 1;
defparam ram_block1a58.port_b_first_address = 0;
defparam ram_block1a58.port_b_first_bit_number = 58;
defparam ram_block1a58.port_b_last_address = 7;
defparam ram_block1a58.port_b_logical_ram_depth = 8;
defparam ram_block1a58.port_b_logical_ram_width = 258;
defparam ram_block1a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a58.port_b_read_enable_clock = "clock1";
defparam ram_block1a58.ram_block_type = "auto";

cycloneive_ram_block ram_block1a57(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[57]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a57_PORTBDATAOUT_bus));
defparam ram_block1a57.clk1_output_clock_enable = "ena1";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a57.operation_mode = "dual_port";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 3;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "none";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 0;
defparam ram_block1a57.port_a_first_bit_number = 57;
defparam ram_block1a57.port_a_last_address = 7;
defparam ram_block1a57.port_a_logical_ram_depth = 8;
defparam ram_block1a57.port_a_logical_ram_width = 258;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a57.port_b_address_clear = "none";
defparam ram_block1a57.port_b_address_clock = "clock1";
defparam ram_block1a57.port_b_address_width = 3;
defparam ram_block1a57.port_b_data_out_clear = "none";
defparam ram_block1a57.port_b_data_out_clock = "clock1";
defparam ram_block1a57.port_b_data_width = 1;
defparam ram_block1a57.port_b_first_address = 0;
defparam ram_block1a57.port_b_first_bit_number = 57;
defparam ram_block1a57.port_b_last_address = 7;
defparam ram_block1a57.port_b_logical_ram_depth = 8;
defparam ram_block1a57.port_b_logical_ram_width = 258;
defparam ram_block1a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a57.port_b_read_enable_clock = "clock1";
defparam ram_block1a57.ram_block_type = "auto";

cycloneive_ram_block ram_block1a56(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[56]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a56_PORTBDATAOUT_bus));
defparam ram_block1a56.clk1_output_clock_enable = "ena1";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a56.operation_mode = "dual_port";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 3;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "none";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 0;
defparam ram_block1a56.port_a_first_bit_number = 56;
defparam ram_block1a56.port_a_last_address = 7;
defparam ram_block1a56.port_a_logical_ram_depth = 8;
defparam ram_block1a56.port_a_logical_ram_width = 258;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a56.port_b_address_clear = "none";
defparam ram_block1a56.port_b_address_clock = "clock1";
defparam ram_block1a56.port_b_address_width = 3;
defparam ram_block1a56.port_b_data_out_clear = "none";
defparam ram_block1a56.port_b_data_out_clock = "clock1";
defparam ram_block1a56.port_b_data_width = 1;
defparam ram_block1a56.port_b_first_address = 0;
defparam ram_block1a56.port_b_first_bit_number = 56;
defparam ram_block1a56.port_b_last_address = 7;
defparam ram_block1a56.port_b_logical_ram_depth = 8;
defparam ram_block1a56.port_b_logical_ram_width = 258;
defparam ram_block1a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a56.port_b_read_enable_clock = "clock1";
defparam ram_block1a56.ram_block_type = "auto";

cycloneive_ram_block ram_block1a55(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[55]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a55_PORTBDATAOUT_bus));
defparam ram_block1a55.clk1_output_clock_enable = "ena1";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a55.operation_mode = "dual_port";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 3;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "none";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 0;
defparam ram_block1a55.port_a_first_bit_number = 55;
defparam ram_block1a55.port_a_last_address = 7;
defparam ram_block1a55.port_a_logical_ram_depth = 8;
defparam ram_block1a55.port_a_logical_ram_width = 258;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a55.port_b_address_clear = "none";
defparam ram_block1a55.port_b_address_clock = "clock1";
defparam ram_block1a55.port_b_address_width = 3;
defparam ram_block1a55.port_b_data_out_clear = "none";
defparam ram_block1a55.port_b_data_out_clock = "clock1";
defparam ram_block1a55.port_b_data_width = 1;
defparam ram_block1a55.port_b_first_address = 0;
defparam ram_block1a55.port_b_first_bit_number = 55;
defparam ram_block1a55.port_b_last_address = 7;
defparam ram_block1a55.port_b_logical_ram_depth = 8;
defparam ram_block1a55.port_b_logical_ram_width = 258;
defparam ram_block1a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a55.port_b_read_enable_clock = "clock1";
defparam ram_block1a55.ram_block_type = "auto";

cycloneive_ram_block ram_block1a54(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[54]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a54_PORTBDATAOUT_bus));
defparam ram_block1a54.clk1_output_clock_enable = "ena1";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a54.operation_mode = "dual_port";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 3;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "none";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 0;
defparam ram_block1a54.port_a_first_bit_number = 54;
defparam ram_block1a54.port_a_last_address = 7;
defparam ram_block1a54.port_a_logical_ram_depth = 8;
defparam ram_block1a54.port_a_logical_ram_width = 258;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a54.port_b_address_clear = "none";
defparam ram_block1a54.port_b_address_clock = "clock1";
defparam ram_block1a54.port_b_address_width = 3;
defparam ram_block1a54.port_b_data_out_clear = "none";
defparam ram_block1a54.port_b_data_out_clock = "clock1";
defparam ram_block1a54.port_b_data_width = 1;
defparam ram_block1a54.port_b_first_address = 0;
defparam ram_block1a54.port_b_first_bit_number = 54;
defparam ram_block1a54.port_b_last_address = 7;
defparam ram_block1a54.port_b_logical_ram_depth = 8;
defparam ram_block1a54.port_b_logical_ram_width = 258;
defparam ram_block1a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a54.port_b_read_enable_clock = "clock1";
defparam ram_block1a54.ram_block_type = "auto";

cycloneive_ram_block ram_block1a53(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[53]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a53_PORTBDATAOUT_bus));
defparam ram_block1a53.clk1_output_clock_enable = "ena1";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a53.operation_mode = "dual_port";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 3;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "none";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 0;
defparam ram_block1a53.port_a_first_bit_number = 53;
defparam ram_block1a53.port_a_last_address = 7;
defparam ram_block1a53.port_a_logical_ram_depth = 8;
defparam ram_block1a53.port_a_logical_ram_width = 258;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a53.port_b_address_clear = "none";
defparam ram_block1a53.port_b_address_clock = "clock1";
defparam ram_block1a53.port_b_address_width = 3;
defparam ram_block1a53.port_b_data_out_clear = "none";
defparam ram_block1a53.port_b_data_out_clock = "clock1";
defparam ram_block1a53.port_b_data_width = 1;
defparam ram_block1a53.port_b_first_address = 0;
defparam ram_block1a53.port_b_first_bit_number = 53;
defparam ram_block1a53.port_b_last_address = 7;
defparam ram_block1a53.port_b_logical_ram_depth = 8;
defparam ram_block1a53.port_b_logical_ram_width = 258;
defparam ram_block1a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a53.port_b_read_enable_clock = "clock1";
defparam ram_block1a53.ram_block_type = "auto";

cycloneive_ram_block ram_block1a52(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[52]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a52_PORTBDATAOUT_bus));
defparam ram_block1a52.clk1_output_clock_enable = "ena1";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a52.operation_mode = "dual_port";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 3;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "none";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 0;
defparam ram_block1a52.port_a_first_bit_number = 52;
defparam ram_block1a52.port_a_last_address = 7;
defparam ram_block1a52.port_a_logical_ram_depth = 8;
defparam ram_block1a52.port_a_logical_ram_width = 258;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a52.port_b_address_clear = "none";
defparam ram_block1a52.port_b_address_clock = "clock1";
defparam ram_block1a52.port_b_address_width = 3;
defparam ram_block1a52.port_b_data_out_clear = "none";
defparam ram_block1a52.port_b_data_out_clock = "clock1";
defparam ram_block1a52.port_b_data_width = 1;
defparam ram_block1a52.port_b_first_address = 0;
defparam ram_block1a52.port_b_first_bit_number = 52;
defparam ram_block1a52.port_b_last_address = 7;
defparam ram_block1a52.port_b_logical_ram_depth = 8;
defparam ram_block1a52.port_b_logical_ram_width = 258;
defparam ram_block1a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a52.port_b_read_enable_clock = "clock1";
defparam ram_block1a52.ram_block_type = "auto";

cycloneive_ram_block ram_block1a90(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[90]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a90_PORTBDATAOUT_bus));
defparam ram_block1a90.clk1_output_clock_enable = "ena1";
defparam ram_block1a90.data_interleave_offset_in_bits = 1;
defparam ram_block1a90.data_interleave_width_in_bits = 1;
defparam ram_block1a90.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a90.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a90.operation_mode = "dual_port";
defparam ram_block1a90.port_a_address_clear = "none";
defparam ram_block1a90.port_a_address_width = 3;
defparam ram_block1a90.port_a_data_out_clear = "none";
defparam ram_block1a90.port_a_data_out_clock = "none";
defparam ram_block1a90.port_a_data_width = 1;
defparam ram_block1a90.port_a_first_address = 0;
defparam ram_block1a90.port_a_first_bit_number = 90;
defparam ram_block1a90.port_a_last_address = 7;
defparam ram_block1a90.port_a_logical_ram_depth = 8;
defparam ram_block1a90.port_a_logical_ram_width = 258;
defparam ram_block1a90.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a90.port_b_address_clear = "none";
defparam ram_block1a90.port_b_address_clock = "clock1";
defparam ram_block1a90.port_b_address_width = 3;
defparam ram_block1a90.port_b_data_out_clear = "none";
defparam ram_block1a90.port_b_data_out_clock = "clock1";
defparam ram_block1a90.port_b_data_width = 1;
defparam ram_block1a90.port_b_first_address = 0;
defparam ram_block1a90.port_b_first_bit_number = 90;
defparam ram_block1a90.port_b_last_address = 7;
defparam ram_block1a90.port_b_logical_ram_depth = 8;
defparam ram_block1a90.port_b_logical_ram_width = 258;
defparam ram_block1a90.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a90.port_b_read_enable_clock = "clock1";
defparam ram_block1a90.ram_block_type = "auto";

cycloneive_ram_block ram_block1a89(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[89]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a89_PORTBDATAOUT_bus));
defparam ram_block1a89.clk1_output_clock_enable = "ena1";
defparam ram_block1a89.data_interleave_offset_in_bits = 1;
defparam ram_block1a89.data_interleave_width_in_bits = 1;
defparam ram_block1a89.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a89.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a89.operation_mode = "dual_port";
defparam ram_block1a89.port_a_address_clear = "none";
defparam ram_block1a89.port_a_address_width = 3;
defparam ram_block1a89.port_a_data_out_clear = "none";
defparam ram_block1a89.port_a_data_out_clock = "none";
defparam ram_block1a89.port_a_data_width = 1;
defparam ram_block1a89.port_a_first_address = 0;
defparam ram_block1a89.port_a_first_bit_number = 89;
defparam ram_block1a89.port_a_last_address = 7;
defparam ram_block1a89.port_a_logical_ram_depth = 8;
defparam ram_block1a89.port_a_logical_ram_width = 258;
defparam ram_block1a89.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a89.port_b_address_clear = "none";
defparam ram_block1a89.port_b_address_clock = "clock1";
defparam ram_block1a89.port_b_address_width = 3;
defparam ram_block1a89.port_b_data_out_clear = "none";
defparam ram_block1a89.port_b_data_out_clock = "clock1";
defparam ram_block1a89.port_b_data_width = 1;
defparam ram_block1a89.port_b_first_address = 0;
defparam ram_block1a89.port_b_first_bit_number = 89;
defparam ram_block1a89.port_b_last_address = 7;
defparam ram_block1a89.port_b_logical_ram_depth = 8;
defparam ram_block1a89.port_b_logical_ram_width = 258;
defparam ram_block1a89.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a89.port_b_read_enable_clock = "clock1";
defparam ram_block1a89.ram_block_type = "auto";

cycloneive_ram_block ram_block1a88(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[88]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a88_PORTBDATAOUT_bus));
defparam ram_block1a88.clk1_output_clock_enable = "ena1";
defparam ram_block1a88.data_interleave_offset_in_bits = 1;
defparam ram_block1a88.data_interleave_width_in_bits = 1;
defparam ram_block1a88.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a88.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a88.operation_mode = "dual_port";
defparam ram_block1a88.port_a_address_clear = "none";
defparam ram_block1a88.port_a_address_width = 3;
defparam ram_block1a88.port_a_data_out_clear = "none";
defparam ram_block1a88.port_a_data_out_clock = "none";
defparam ram_block1a88.port_a_data_width = 1;
defparam ram_block1a88.port_a_first_address = 0;
defparam ram_block1a88.port_a_first_bit_number = 88;
defparam ram_block1a88.port_a_last_address = 7;
defparam ram_block1a88.port_a_logical_ram_depth = 8;
defparam ram_block1a88.port_a_logical_ram_width = 258;
defparam ram_block1a88.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a88.port_b_address_clear = "none";
defparam ram_block1a88.port_b_address_clock = "clock1";
defparam ram_block1a88.port_b_address_width = 3;
defparam ram_block1a88.port_b_data_out_clear = "none";
defparam ram_block1a88.port_b_data_out_clock = "clock1";
defparam ram_block1a88.port_b_data_width = 1;
defparam ram_block1a88.port_b_first_address = 0;
defparam ram_block1a88.port_b_first_bit_number = 88;
defparam ram_block1a88.port_b_last_address = 7;
defparam ram_block1a88.port_b_logical_ram_depth = 8;
defparam ram_block1a88.port_b_logical_ram_width = 258;
defparam ram_block1a88.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a88.port_b_read_enable_clock = "clock1";
defparam ram_block1a88.ram_block_type = "auto";

cycloneive_ram_block ram_block1a87(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[87]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a87_PORTBDATAOUT_bus));
defparam ram_block1a87.clk1_output_clock_enable = "ena1";
defparam ram_block1a87.data_interleave_offset_in_bits = 1;
defparam ram_block1a87.data_interleave_width_in_bits = 1;
defparam ram_block1a87.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a87.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a87.operation_mode = "dual_port";
defparam ram_block1a87.port_a_address_clear = "none";
defparam ram_block1a87.port_a_address_width = 3;
defparam ram_block1a87.port_a_data_out_clear = "none";
defparam ram_block1a87.port_a_data_out_clock = "none";
defparam ram_block1a87.port_a_data_width = 1;
defparam ram_block1a87.port_a_first_address = 0;
defparam ram_block1a87.port_a_first_bit_number = 87;
defparam ram_block1a87.port_a_last_address = 7;
defparam ram_block1a87.port_a_logical_ram_depth = 8;
defparam ram_block1a87.port_a_logical_ram_width = 258;
defparam ram_block1a87.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a87.port_b_address_clear = "none";
defparam ram_block1a87.port_b_address_clock = "clock1";
defparam ram_block1a87.port_b_address_width = 3;
defparam ram_block1a87.port_b_data_out_clear = "none";
defparam ram_block1a87.port_b_data_out_clock = "clock1";
defparam ram_block1a87.port_b_data_width = 1;
defparam ram_block1a87.port_b_first_address = 0;
defparam ram_block1a87.port_b_first_bit_number = 87;
defparam ram_block1a87.port_b_last_address = 7;
defparam ram_block1a87.port_b_logical_ram_depth = 8;
defparam ram_block1a87.port_b_logical_ram_width = 258;
defparam ram_block1a87.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a87.port_b_read_enable_clock = "clock1";
defparam ram_block1a87.ram_block_type = "auto";

cycloneive_ram_block ram_block1a86(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[86]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a86_PORTBDATAOUT_bus));
defparam ram_block1a86.clk1_output_clock_enable = "ena1";
defparam ram_block1a86.data_interleave_offset_in_bits = 1;
defparam ram_block1a86.data_interleave_width_in_bits = 1;
defparam ram_block1a86.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a86.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a86.operation_mode = "dual_port";
defparam ram_block1a86.port_a_address_clear = "none";
defparam ram_block1a86.port_a_address_width = 3;
defparam ram_block1a86.port_a_data_out_clear = "none";
defparam ram_block1a86.port_a_data_out_clock = "none";
defparam ram_block1a86.port_a_data_width = 1;
defparam ram_block1a86.port_a_first_address = 0;
defparam ram_block1a86.port_a_first_bit_number = 86;
defparam ram_block1a86.port_a_last_address = 7;
defparam ram_block1a86.port_a_logical_ram_depth = 8;
defparam ram_block1a86.port_a_logical_ram_width = 258;
defparam ram_block1a86.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a86.port_b_address_clear = "none";
defparam ram_block1a86.port_b_address_clock = "clock1";
defparam ram_block1a86.port_b_address_width = 3;
defparam ram_block1a86.port_b_data_out_clear = "none";
defparam ram_block1a86.port_b_data_out_clock = "clock1";
defparam ram_block1a86.port_b_data_width = 1;
defparam ram_block1a86.port_b_first_address = 0;
defparam ram_block1a86.port_b_first_bit_number = 86;
defparam ram_block1a86.port_b_last_address = 7;
defparam ram_block1a86.port_b_logical_ram_depth = 8;
defparam ram_block1a86.port_b_logical_ram_width = 258;
defparam ram_block1a86.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a86.port_b_read_enable_clock = "clock1";
defparam ram_block1a86.ram_block_type = "auto";

cycloneive_ram_block ram_block1a85(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[85]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a85_PORTBDATAOUT_bus));
defparam ram_block1a85.clk1_output_clock_enable = "ena1";
defparam ram_block1a85.data_interleave_offset_in_bits = 1;
defparam ram_block1a85.data_interleave_width_in_bits = 1;
defparam ram_block1a85.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a85.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a85.operation_mode = "dual_port";
defparam ram_block1a85.port_a_address_clear = "none";
defparam ram_block1a85.port_a_address_width = 3;
defparam ram_block1a85.port_a_data_out_clear = "none";
defparam ram_block1a85.port_a_data_out_clock = "none";
defparam ram_block1a85.port_a_data_width = 1;
defparam ram_block1a85.port_a_first_address = 0;
defparam ram_block1a85.port_a_first_bit_number = 85;
defparam ram_block1a85.port_a_last_address = 7;
defparam ram_block1a85.port_a_logical_ram_depth = 8;
defparam ram_block1a85.port_a_logical_ram_width = 258;
defparam ram_block1a85.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a85.port_b_address_clear = "none";
defparam ram_block1a85.port_b_address_clock = "clock1";
defparam ram_block1a85.port_b_address_width = 3;
defparam ram_block1a85.port_b_data_out_clear = "none";
defparam ram_block1a85.port_b_data_out_clock = "clock1";
defparam ram_block1a85.port_b_data_width = 1;
defparam ram_block1a85.port_b_first_address = 0;
defparam ram_block1a85.port_b_first_bit_number = 85;
defparam ram_block1a85.port_b_last_address = 7;
defparam ram_block1a85.port_b_logical_ram_depth = 8;
defparam ram_block1a85.port_b_logical_ram_width = 258;
defparam ram_block1a85.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a85.port_b_read_enable_clock = "clock1";
defparam ram_block1a85.ram_block_type = "auto";

cycloneive_ram_block ram_block1a84(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[84]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a84_PORTBDATAOUT_bus));
defparam ram_block1a84.clk1_output_clock_enable = "ena1";
defparam ram_block1a84.data_interleave_offset_in_bits = 1;
defparam ram_block1a84.data_interleave_width_in_bits = 1;
defparam ram_block1a84.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a84.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a84.operation_mode = "dual_port";
defparam ram_block1a84.port_a_address_clear = "none";
defparam ram_block1a84.port_a_address_width = 3;
defparam ram_block1a84.port_a_data_out_clear = "none";
defparam ram_block1a84.port_a_data_out_clock = "none";
defparam ram_block1a84.port_a_data_width = 1;
defparam ram_block1a84.port_a_first_address = 0;
defparam ram_block1a84.port_a_first_bit_number = 84;
defparam ram_block1a84.port_a_last_address = 7;
defparam ram_block1a84.port_a_logical_ram_depth = 8;
defparam ram_block1a84.port_a_logical_ram_width = 258;
defparam ram_block1a84.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a84.port_b_address_clear = "none";
defparam ram_block1a84.port_b_address_clock = "clock1";
defparam ram_block1a84.port_b_address_width = 3;
defparam ram_block1a84.port_b_data_out_clear = "none";
defparam ram_block1a84.port_b_data_out_clock = "clock1";
defparam ram_block1a84.port_b_data_width = 1;
defparam ram_block1a84.port_b_first_address = 0;
defparam ram_block1a84.port_b_first_bit_number = 84;
defparam ram_block1a84.port_b_last_address = 7;
defparam ram_block1a84.port_b_logical_ram_depth = 8;
defparam ram_block1a84.port_b_logical_ram_width = 258;
defparam ram_block1a84.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a84.port_b_read_enable_clock = "clock1";
defparam ram_block1a84.ram_block_type = "auto";

cycloneive_ram_block ram_block1a154(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[154]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a154_PORTBDATAOUT_bus));
defparam ram_block1a154.clk1_output_clock_enable = "ena1";
defparam ram_block1a154.data_interleave_offset_in_bits = 1;
defparam ram_block1a154.data_interleave_width_in_bits = 1;
defparam ram_block1a154.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a154.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a154.operation_mode = "dual_port";
defparam ram_block1a154.port_a_address_clear = "none";
defparam ram_block1a154.port_a_address_width = 3;
defparam ram_block1a154.port_a_data_out_clear = "none";
defparam ram_block1a154.port_a_data_out_clock = "none";
defparam ram_block1a154.port_a_data_width = 1;
defparam ram_block1a154.port_a_first_address = 0;
defparam ram_block1a154.port_a_first_bit_number = 154;
defparam ram_block1a154.port_a_last_address = 7;
defparam ram_block1a154.port_a_logical_ram_depth = 8;
defparam ram_block1a154.port_a_logical_ram_width = 258;
defparam ram_block1a154.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a154.port_b_address_clear = "none";
defparam ram_block1a154.port_b_address_clock = "clock1";
defparam ram_block1a154.port_b_address_width = 3;
defparam ram_block1a154.port_b_data_out_clear = "none";
defparam ram_block1a154.port_b_data_out_clock = "clock1";
defparam ram_block1a154.port_b_data_width = 1;
defparam ram_block1a154.port_b_first_address = 0;
defparam ram_block1a154.port_b_first_bit_number = 154;
defparam ram_block1a154.port_b_last_address = 7;
defparam ram_block1a154.port_b_logical_ram_depth = 8;
defparam ram_block1a154.port_b_logical_ram_width = 258;
defparam ram_block1a154.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a154.port_b_read_enable_clock = "clock1";
defparam ram_block1a154.ram_block_type = "auto";

cycloneive_ram_block ram_block1a153(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[153]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a153_PORTBDATAOUT_bus));
defparam ram_block1a153.clk1_output_clock_enable = "ena1";
defparam ram_block1a153.data_interleave_offset_in_bits = 1;
defparam ram_block1a153.data_interleave_width_in_bits = 1;
defparam ram_block1a153.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a153.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a153.operation_mode = "dual_port";
defparam ram_block1a153.port_a_address_clear = "none";
defparam ram_block1a153.port_a_address_width = 3;
defparam ram_block1a153.port_a_data_out_clear = "none";
defparam ram_block1a153.port_a_data_out_clock = "none";
defparam ram_block1a153.port_a_data_width = 1;
defparam ram_block1a153.port_a_first_address = 0;
defparam ram_block1a153.port_a_first_bit_number = 153;
defparam ram_block1a153.port_a_last_address = 7;
defparam ram_block1a153.port_a_logical_ram_depth = 8;
defparam ram_block1a153.port_a_logical_ram_width = 258;
defparam ram_block1a153.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a153.port_b_address_clear = "none";
defparam ram_block1a153.port_b_address_clock = "clock1";
defparam ram_block1a153.port_b_address_width = 3;
defparam ram_block1a153.port_b_data_out_clear = "none";
defparam ram_block1a153.port_b_data_out_clock = "clock1";
defparam ram_block1a153.port_b_data_width = 1;
defparam ram_block1a153.port_b_first_address = 0;
defparam ram_block1a153.port_b_first_bit_number = 153;
defparam ram_block1a153.port_b_last_address = 7;
defparam ram_block1a153.port_b_logical_ram_depth = 8;
defparam ram_block1a153.port_b_logical_ram_width = 258;
defparam ram_block1a153.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a153.port_b_read_enable_clock = "clock1";
defparam ram_block1a153.ram_block_type = "auto";

cycloneive_ram_block ram_block1a152(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[152]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a152_PORTBDATAOUT_bus));
defparam ram_block1a152.clk1_output_clock_enable = "ena1";
defparam ram_block1a152.data_interleave_offset_in_bits = 1;
defparam ram_block1a152.data_interleave_width_in_bits = 1;
defparam ram_block1a152.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a152.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a152.operation_mode = "dual_port";
defparam ram_block1a152.port_a_address_clear = "none";
defparam ram_block1a152.port_a_address_width = 3;
defparam ram_block1a152.port_a_data_out_clear = "none";
defparam ram_block1a152.port_a_data_out_clock = "none";
defparam ram_block1a152.port_a_data_width = 1;
defparam ram_block1a152.port_a_first_address = 0;
defparam ram_block1a152.port_a_first_bit_number = 152;
defparam ram_block1a152.port_a_last_address = 7;
defparam ram_block1a152.port_a_logical_ram_depth = 8;
defparam ram_block1a152.port_a_logical_ram_width = 258;
defparam ram_block1a152.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a152.port_b_address_clear = "none";
defparam ram_block1a152.port_b_address_clock = "clock1";
defparam ram_block1a152.port_b_address_width = 3;
defparam ram_block1a152.port_b_data_out_clear = "none";
defparam ram_block1a152.port_b_data_out_clock = "clock1";
defparam ram_block1a152.port_b_data_width = 1;
defparam ram_block1a152.port_b_first_address = 0;
defparam ram_block1a152.port_b_first_bit_number = 152;
defparam ram_block1a152.port_b_last_address = 7;
defparam ram_block1a152.port_b_logical_ram_depth = 8;
defparam ram_block1a152.port_b_logical_ram_width = 258;
defparam ram_block1a152.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a152.port_b_read_enable_clock = "clock1";
defparam ram_block1a152.ram_block_type = "auto";

cycloneive_ram_block ram_block1a151(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[151]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a151_PORTBDATAOUT_bus));
defparam ram_block1a151.clk1_output_clock_enable = "ena1";
defparam ram_block1a151.data_interleave_offset_in_bits = 1;
defparam ram_block1a151.data_interleave_width_in_bits = 1;
defparam ram_block1a151.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a151.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a151.operation_mode = "dual_port";
defparam ram_block1a151.port_a_address_clear = "none";
defparam ram_block1a151.port_a_address_width = 3;
defparam ram_block1a151.port_a_data_out_clear = "none";
defparam ram_block1a151.port_a_data_out_clock = "none";
defparam ram_block1a151.port_a_data_width = 1;
defparam ram_block1a151.port_a_first_address = 0;
defparam ram_block1a151.port_a_first_bit_number = 151;
defparam ram_block1a151.port_a_last_address = 7;
defparam ram_block1a151.port_a_logical_ram_depth = 8;
defparam ram_block1a151.port_a_logical_ram_width = 258;
defparam ram_block1a151.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a151.port_b_address_clear = "none";
defparam ram_block1a151.port_b_address_clock = "clock1";
defparam ram_block1a151.port_b_address_width = 3;
defparam ram_block1a151.port_b_data_out_clear = "none";
defparam ram_block1a151.port_b_data_out_clock = "clock1";
defparam ram_block1a151.port_b_data_width = 1;
defparam ram_block1a151.port_b_first_address = 0;
defparam ram_block1a151.port_b_first_bit_number = 151;
defparam ram_block1a151.port_b_last_address = 7;
defparam ram_block1a151.port_b_logical_ram_depth = 8;
defparam ram_block1a151.port_b_logical_ram_width = 258;
defparam ram_block1a151.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a151.port_b_read_enable_clock = "clock1";
defparam ram_block1a151.ram_block_type = "auto";

cycloneive_ram_block ram_block1a150(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[150]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a150_PORTBDATAOUT_bus));
defparam ram_block1a150.clk1_output_clock_enable = "ena1";
defparam ram_block1a150.data_interleave_offset_in_bits = 1;
defparam ram_block1a150.data_interleave_width_in_bits = 1;
defparam ram_block1a150.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a150.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a150.operation_mode = "dual_port";
defparam ram_block1a150.port_a_address_clear = "none";
defparam ram_block1a150.port_a_address_width = 3;
defparam ram_block1a150.port_a_data_out_clear = "none";
defparam ram_block1a150.port_a_data_out_clock = "none";
defparam ram_block1a150.port_a_data_width = 1;
defparam ram_block1a150.port_a_first_address = 0;
defparam ram_block1a150.port_a_first_bit_number = 150;
defparam ram_block1a150.port_a_last_address = 7;
defparam ram_block1a150.port_a_logical_ram_depth = 8;
defparam ram_block1a150.port_a_logical_ram_width = 258;
defparam ram_block1a150.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a150.port_b_address_clear = "none";
defparam ram_block1a150.port_b_address_clock = "clock1";
defparam ram_block1a150.port_b_address_width = 3;
defparam ram_block1a150.port_b_data_out_clear = "none";
defparam ram_block1a150.port_b_data_out_clock = "clock1";
defparam ram_block1a150.port_b_data_width = 1;
defparam ram_block1a150.port_b_first_address = 0;
defparam ram_block1a150.port_b_first_bit_number = 150;
defparam ram_block1a150.port_b_last_address = 7;
defparam ram_block1a150.port_b_logical_ram_depth = 8;
defparam ram_block1a150.port_b_logical_ram_width = 258;
defparam ram_block1a150.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a150.port_b_read_enable_clock = "clock1";
defparam ram_block1a150.ram_block_type = "auto";

cycloneive_ram_block ram_block1a149(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[149]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a149_PORTBDATAOUT_bus));
defparam ram_block1a149.clk1_output_clock_enable = "ena1";
defparam ram_block1a149.data_interleave_offset_in_bits = 1;
defparam ram_block1a149.data_interleave_width_in_bits = 1;
defparam ram_block1a149.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a149.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a149.operation_mode = "dual_port";
defparam ram_block1a149.port_a_address_clear = "none";
defparam ram_block1a149.port_a_address_width = 3;
defparam ram_block1a149.port_a_data_out_clear = "none";
defparam ram_block1a149.port_a_data_out_clock = "none";
defparam ram_block1a149.port_a_data_width = 1;
defparam ram_block1a149.port_a_first_address = 0;
defparam ram_block1a149.port_a_first_bit_number = 149;
defparam ram_block1a149.port_a_last_address = 7;
defparam ram_block1a149.port_a_logical_ram_depth = 8;
defparam ram_block1a149.port_a_logical_ram_width = 258;
defparam ram_block1a149.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a149.port_b_address_clear = "none";
defparam ram_block1a149.port_b_address_clock = "clock1";
defparam ram_block1a149.port_b_address_width = 3;
defparam ram_block1a149.port_b_data_out_clear = "none";
defparam ram_block1a149.port_b_data_out_clock = "clock1";
defparam ram_block1a149.port_b_data_width = 1;
defparam ram_block1a149.port_b_first_address = 0;
defparam ram_block1a149.port_b_first_bit_number = 149;
defparam ram_block1a149.port_b_last_address = 7;
defparam ram_block1a149.port_b_logical_ram_depth = 8;
defparam ram_block1a149.port_b_logical_ram_width = 258;
defparam ram_block1a149.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a149.port_b_read_enable_clock = "clock1";
defparam ram_block1a149.ram_block_type = "auto";

cycloneive_ram_block ram_block1a148(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[148]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a148_PORTBDATAOUT_bus));
defparam ram_block1a148.clk1_output_clock_enable = "ena1";
defparam ram_block1a148.data_interleave_offset_in_bits = 1;
defparam ram_block1a148.data_interleave_width_in_bits = 1;
defparam ram_block1a148.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a148.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a148.operation_mode = "dual_port";
defparam ram_block1a148.port_a_address_clear = "none";
defparam ram_block1a148.port_a_address_width = 3;
defparam ram_block1a148.port_a_data_out_clear = "none";
defparam ram_block1a148.port_a_data_out_clock = "none";
defparam ram_block1a148.port_a_data_width = 1;
defparam ram_block1a148.port_a_first_address = 0;
defparam ram_block1a148.port_a_first_bit_number = 148;
defparam ram_block1a148.port_a_last_address = 7;
defparam ram_block1a148.port_a_logical_ram_depth = 8;
defparam ram_block1a148.port_a_logical_ram_width = 258;
defparam ram_block1a148.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a148.port_b_address_clear = "none";
defparam ram_block1a148.port_b_address_clock = "clock1";
defparam ram_block1a148.port_b_address_width = 3;
defparam ram_block1a148.port_b_data_out_clear = "none";
defparam ram_block1a148.port_b_data_out_clock = "clock1";
defparam ram_block1a148.port_b_data_width = 1;
defparam ram_block1a148.port_b_first_address = 0;
defparam ram_block1a148.port_b_first_bit_number = 148;
defparam ram_block1a148.port_b_last_address = 7;
defparam ram_block1a148.port_b_logical_ram_depth = 8;
defparam ram_block1a148.port_b_logical_ram_width = 258;
defparam ram_block1a148.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a148.port_b_read_enable_clock = "clock1";
defparam ram_block1a148.ram_block_type = "auto";

cycloneive_ram_block ram_block1a218(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[218]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a218_PORTBDATAOUT_bus));
defparam ram_block1a218.clk1_output_clock_enable = "ena1";
defparam ram_block1a218.data_interleave_offset_in_bits = 1;
defparam ram_block1a218.data_interleave_width_in_bits = 1;
defparam ram_block1a218.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a218.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a218.operation_mode = "dual_port";
defparam ram_block1a218.port_a_address_clear = "none";
defparam ram_block1a218.port_a_address_width = 3;
defparam ram_block1a218.port_a_data_out_clear = "none";
defparam ram_block1a218.port_a_data_out_clock = "none";
defparam ram_block1a218.port_a_data_width = 1;
defparam ram_block1a218.port_a_first_address = 0;
defparam ram_block1a218.port_a_first_bit_number = 218;
defparam ram_block1a218.port_a_last_address = 7;
defparam ram_block1a218.port_a_logical_ram_depth = 8;
defparam ram_block1a218.port_a_logical_ram_width = 258;
defparam ram_block1a218.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a218.port_b_address_clear = "none";
defparam ram_block1a218.port_b_address_clock = "clock1";
defparam ram_block1a218.port_b_address_width = 3;
defparam ram_block1a218.port_b_data_out_clear = "none";
defparam ram_block1a218.port_b_data_out_clock = "clock1";
defparam ram_block1a218.port_b_data_width = 1;
defparam ram_block1a218.port_b_first_address = 0;
defparam ram_block1a218.port_b_first_bit_number = 218;
defparam ram_block1a218.port_b_last_address = 7;
defparam ram_block1a218.port_b_logical_ram_depth = 8;
defparam ram_block1a218.port_b_logical_ram_width = 258;
defparam ram_block1a218.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a218.port_b_read_enable_clock = "clock1";
defparam ram_block1a218.ram_block_type = "auto";

cycloneive_ram_block ram_block1a217(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[217]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a217_PORTBDATAOUT_bus));
defparam ram_block1a217.clk1_output_clock_enable = "ena1";
defparam ram_block1a217.data_interleave_offset_in_bits = 1;
defparam ram_block1a217.data_interleave_width_in_bits = 1;
defparam ram_block1a217.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a217.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a217.operation_mode = "dual_port";
defparam ram_block1a217.port_a_address_clear = "none";
defparam ram_block1a217.port_a_address_width = 3;
defparam ram_block1a217.port_a_data_out_clear = "none";
defparam ram_block1a217.port_a_data_out_clock = "none";
defparam ram_block1a217.port_a_data_width = 1;
defparam ram_block1a217.port_a_first_address = 0;
defparam ram_block1a217.port_a_first_bit_number = 217;
defparam ram_block1a217.port_a_last_address = 7;
defparam ram_block1a217.port_a_logical_ram_depth = 8;
defparam ram_block1a217.port_a_logical_ram_width = 258;
defparam ram_block1a217.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a217.port_b_address_clear = "none";
defparam ram_block1a217.port_b_address_clock = "clock1";
defparam ram_block1a217.port_b_address_width = 3;
defparam ram_block1a217.port_b_data_out_clear = "none";
defparam ram_block1a217.port_b_data_out_clock = "clock1";
defparam ram_block1a217.port_b_data_width = 1;
defparam ram_block1a217.port_b_first_address = 0;
defparam ram_block1a217.port_b_first_bit_number = 217;
defparam ram_block1a217.port_b_last_address = 7;
defparam ram_block1a217.port_b_logical_ram_depth = 8;
defparam ram_block1a217.port_b_logical_ram_width = 258;
defparam ram_block1a217.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a217.port_b_read_enable_clock = "clock1";
defparam ram_block1a217.ram_block_type = "auto";

cycloneive_ram_block ram_block1a216(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[216]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a216_PORTBDATAOUT_bus));
defparam ram_block1a216.clk1_output_clock_enable = "ena1";
defparam ram_block1a216.data_interleave_offset_in_bits = 1;
defparam ram_block1a216.data_interleave_width_in_bits = 1;
defparam ram_block1a216.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a216.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a216.operation_mode = "dual_port";
defparam ram_block1a216.port_a_address_clear = "none";
defparam ram_block1a216.port_a_address_width = 3;
defparam ram_block1a216.port_a_data_out_clear = "none";
defparam ram_block1a216.port_a_data_out_clock = "none";
defparam ram_block1a216.port_a_data_width = 1;
defparam ram_block1a216.port_a_first_address = 0;
defparam ram_block1a216.port_a_first_bit_number = 216;
defparam ram_block1a216.port_a_last_address = 7;
defparam ram_block1a216.port_a_logical_ram_depth = 8;
defparam ram_block1a216.port_a_logical_ram_width = 258;
defparam ram_block1a216.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a216.port_b_address_clear = "none";
defparam ram_block1a216.port_b_address_clock = "clock1";
defparam ram_block1a216.port_b_address_width = 3;
defparam ram_block1a216.port_b_data_out_clear = "none";
defparam ram_block1a216.port_b_data_out_clock = "clock1";
defparam ram_block1a216.port_b_data_width = 1;
defparam ram_block1a216.port_b_first_address = 0;
defparam ram_block1a216.port_b_first_bit_number = 216;
defparam ram_block1a216.port_b_last_address = 7;
defparam ram_block1a216.port_b_logical_ram_depth = 8;
defparam ram_block1a216.port_b_logical_ram_width = 258;
defparam ram_block1a216.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a216.port_b_read_enable_clock = "clock1";
defparam ram_block1a216.ram_block_type = "auto";

cycloneive_ram_block ram_block1a215(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[215]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a215_PORTBDATAOUT_bus));
defparam ram_block1a215.clk1_output_clock_enable = "ena1";
defparam ram_block1a215.data_interleave_offset_in_bits = 1;
defparam ram_block1a215.data_interleave_width_in_bits = 1;
defparam ram_block1a215.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a215.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a215.operation_mode = "dual_port";
defparam ram_block1a215.port_a_address_clear = "none";
defparam ram_block1a215.port_a_address_width = 3;
defparam ram_block1a215.port_a_data_out_clear = "none";
defparam ram_block1a215.port_a_data_out_clock = "none";
defparam ram_block1a215.port_a_data_width = 1;
defparam ram_block1a215.port_a_first_address = 0;
defparam ram_block1a215.port_a_first_bit_number = 215;
defparam ram_block1a215.port_a_last_address = 7;
defparam ram_block1a215.port_a_logical_ram_depth = 8;
defparam ram_block1a215.port_a_logical_ram_width = 258;
defparam ram_block1a215.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a215.port_b_address_clear = "none";
defparam ram_block1a215.port_b_address_clock = "clock1";
defparam ram_block1a215.port_b_address_width = 3;
defparam ram_block1a215.port_b_data_out_clear = "none";
defparam ram_block1a215.port_b_data_out_clock = "clock1";
defparam ram_block1a215.port_b_data_width = 1;
defparam ram_block1a215.port_b_first_address = 0;
defparam ram_block1a215.port_b_first_bit_number = 215;
defparam ram_block1a215.port_b_last_address = 7;
defparam ram_block1a215.port_b_logical_ram_depth = 8;
defparam ram_block1a215.port_b_logical_ram_width = 258;
defparam ram_block1a215.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a215.port_b_read_enable_clock = "clock1";
defparam ram_block1a215.ram_block_type = "auto";

cycloneive_ram_block ram_block1a214(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[214]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a214_PORTBDATAOUT_bus));
defparam ram_block1a214.clk1_output_clock_enable = "ena1";
defparam ram_block1a214.data_interleave_offset_in_bits = 1;
defparam ram_block1a214.data_interleave_width_in_bits = 1;
defparam ram_block1a214.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a214.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a214.operation_mode = "dual_port";
defparam ram_block1a214.port_a_address_clear = "none";
defparam ram_block1a214.port_a_address_width = 3;
defparam ram_block1a214.port_a_data_out_clear = "none";
defparam ram_block1a214.port_a_data_out_clock = "none";
defparam ram_block1a214.port_a_data_width = 1;
defparam ram_block1a214.port_a_first_address = 0;
defparam ram_block1a214.port_a_first_bit_number = 214;
defparam ram_block1a214.port_a_last_address = 7;
defparam ram_block1a214.port_a_logical_ram_depth = 8;
defparam ram_block1a214.port_a_logical_ram_width = 258;
defparam ram_block1a214.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a214.port_b_address_clear = "none";
defparam ram_block1a214.port_b_address_clock = "clock1";
defparam ram_block1a214.port_b_address_width = 3;
defparam ram_block1a214.port_b_data_out_clear = "none";
defparam ram_block1a214.port_b_data_out_clock = "clock1";
defparam ram_block1a214.port_b_data_width = 1;
defparam ram_block1a214.port_b_first_address = 0;
defparam ram_block1a214.port_b_first_bit_number = 214;
defparam ram_block1a214.port_b_last_address = 7;
defparam ram_block1a214.port_b_logical_ram_depth = 8;
defparam ram_block1a214.port_b_logical_ram_width = 258;
defparam ram_block1a214.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a214.port_b_read_enable_clock = "clock1";
defparam ram_block1a214.ram_block_type = "auto";

cycloneive_ram_block ram_block1a213(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[213]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a213_PORTBDATAOUT_bus));
defparam ram_block1a213.clk1_output_clock_enable = "ena1";
defparam ram_block1a213.data_interleave_offset_in_bits = 1;
defparam ram_block1a213.data_interleave_width_in_bits = 1;
defparam ram_block1a213.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a213.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a213.operation_mode = "dual_port";
defparam ram_block1a213.port_a_address_clear = "none";
defparam ram_block1a213.port_a_address_width = 3;
defparam ram_block1a213.port_a_data_out_clear = "none";
defparam ram_block1a213.port_a_data_out_clock = "none";
defparam ram_block1a213.port_a_data_width = 1;
defparam ram_block1a213.port_a_first_address = 0;
defparam ram_block1a213.port_a_first_bit_number = 213;
defparam ram_block1a213.port_a_last_address = 7;
defparam ram_block1a213.port_a_logical_ram_depth = 8;
defparam ram_block1a213.port_a_logical_ram_width = 258;
defparam ram_block1a213.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a213.port_b_address_clear = "none";
defparam ram_block1a213.port_b_address_clock = "clock1";
defparam ram_block1a213.port_b_address_width = 3;
defparam ram_block1a213.port_b_data_out_clear = "none";
defparam ram_block1a213.port_b_data_out_clock = "clock1";
defparam ram_block1a213.port_b_data_width = 1;
defparam ram_block1a213.port_b_first_address = 0;
defparam ram_block1a213.port_b_first_bit_number = 213;
defparam ram_block1a213.port_b_last_address = 7;
defparam ram_block1a213.port_b_logical_ram_depth = 8;
defparam ram_block1a213.port_b_logical_ram_width = 258;
defparam ram_block1a213.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a213.port_b_read_enable_clock = "clock1";
defparam ram_block1a213.ram_block_type = "auto";

cycloneive_ram_block ram_block1a212(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[212]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a212_PORTBDATAOUT_bus));
defparam ram_block1a212.clk1_output_clock_enable = "ena1";
defparam ram_block1a212.data_interleave_offset_in_bits = 1;
defparam ram_block1a212.data_interleave_width_in_bits = 1;
defparam ram_block1a212.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a212.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a212.operation_mode = "dual_port";
defparam ram_block1a212.port_a_address_clear = "none";
defparam ram_block1a212.port_a_address_width = 3;
defparam ram_block1a212.port_a_data_out_clear = "none";
defparam ram_block1a212.port_a_data_out_clock = "none";
defparam ram_block1a212.port_a_data_width = 1;
defparam ram_block1a212.port_a_first_address = 0;
defparam ram_block1a212.port_a_first_bit_number = 212;
defparam ram_block1a212.port_a_last_address = 7;
defparam ram_block1a212.port_a_logical_ram_depth = 8;
defparam ram_block1a212.port_a_logical_ram_width = 258;
defparam ram_block1a212.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a212.port_b_address_clear = "none";
defparam ram_block1a212.port_b_address_clock = "clock1";
defparam ram_block1a212.port_b_address_width = 3;
defparam ram_block1a212.port_b_data_out_clear = "none";
defparam ram_block1a212.port_b_data_out_clock = "clock1";
defparam ram_block1a212.port_b_data_width = 1;
defparam ram_block1a212.port_b_first_address = 0;
defparam ram_block1a212.port_b_first_bit_number = 212;
defparam ram_block1a212.port_b_last_address = 7;
defparam ram_block1a212.port_b_logical_ram_depth = 8;
defparam ram_block1a212.port_b_logical_ram_width = 258;
defparam ram_block1a212.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a212.port_b_read_enable_clock = "clock1";
defparam ram_block1a212.ram_block_type = "auto";

cycloneive_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk1_output_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 3;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 7;
defparam ram_block1a26.port_a_logical_ram_depth = 8;
defparam ram_block1a26.port_a_logical_ram_width = 258;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 3;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock1";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 7;
defparam ram_block1a26.port_b_logical_ram_depth = 8;
defparam ram_block1a26.port_b_logical_ram_width = 258;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cycloneive_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk1_output_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 3;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 7;
defparam ram_block1a25.port_a_logical_ram_depth = 8;
defparam ram_block1a25.port_a_logical_ram_width = 258;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 3;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock1";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 7;
defparam ram_block1a25.port_b_logical_ram_depth = 8;
defparam ram_block1a25.port_b_logical_ram_width = 258;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cycloneive_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk1_output_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 3;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 7;
defparam ram_block1a24.port_a_logical_ram_depth = 8;
defparam ram_block1a24.port_a_logical_ram_width = 258;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 3;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock1";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 7;
defparam ram_block1a24.port_b_logical_ram_depth = 8;
defparam ram_block1a24.port_b_logical_ram_width = 258;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cycloneive_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk1_output_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 3;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 7;
defparam ram_block1a23.port_a_logical_ram_depth = 8;
defparam ram_block1a23.port_a_logical_ram_width = 258;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 3;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock1";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 7;
defparam ram_block1a23.port_b_logical_ram_depth = 8;
defparam ram_block1a23.port_b_logical_ram_width = 258;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cycloneive_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk1_output_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 3;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 7;
defparam ram_block1a22.port_a_logical_ram_depth = 8;
defparam ram_block1a22.port_a_logical_ram_width = 258;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 3;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 7;
defparam ram_block1a22.port_b_logical_ram_depth = 8;
defparam ram_block1a22.port_b_logical_ram_width = 258;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cycloneive_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 3;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 7;
defparam ram_block1a21.port_a_logical_ram_depth = 8;
defparam ram_block1a21.port_a_logical_ram_width = 258;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 3;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 7;
defparam ram_block1a21.port_b_logical_ram_depth = 8;
defparam ram_block1a21.port_b_logical_ram_width = 258;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cycloneive_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 3;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 7;
defparam ram_block1a20.port_a_logical_ram_depth = 8;
defparam ram_block1a20.port_a_logical_ram_width = 258;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 3;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 7;
defparam ram_block1a20.port_b_logical_ram_depth = 8;
defparam ram_block1a20.port_b_logical_ram_width = 258;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cycloneive_ram_block ram_block1a74(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[74]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a74_PORTBDATAOUT_bus));
defparam ram_block1a74.clk1_output_clock_enable = "ena1";
defparam ram_block1a74.data_interleave_offset_in_bits = 1;
defparam ram_block1a74.data_interleave_width_in_bits = 1;
defparam ram_block1a74.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a74.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a74.operation_mode = "dual_port";
defparam ram_block1a74.port_a_address_clear = "none";
defparam ram_block1a74.port_a_address_width = 3;
defparam ram_block1a74.port_a_data_out_clear = "none";
defparam ram_block1a74.port_a_data_out_clock = "none";
defparam ram_block1a74.port_a_data_width = 1;
defparam ram_block1a74.port_a_first_address = 0;
defparam ram_block1a74.port_a_first_bit_number = 74;
defparam ram_block1a74.port_a_last_address = 7;
defparam ram_block1a74.port_a_logical_ram_depth = 8;
defparam ram_block1a74.port_a_logical_ram_width = 258;
defparam ram_block1a74.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a74.port_b_address_clear = "none";
defparam ram_block1a74.port_b_address_clock = "clock1";
defparam ram_block1a74.port_b_address_width = 3;
defparam ram_block1a74.port_b_data_out_clear = "none";
defparam ram_block1a74.port_b_data_out_clock = "clock1";
defparam ram_block1a74.port_b_data_width = 1;
defparam ram_block1a74.port_b_first_address = 0;
defparam ram_block1a74.port_b_first_bit_number = 74;
defparam ram_block1a74.port_b_last_address = 7;
defparam ram_block1a74.port_b_logical_ram_depth = 8;
defparam ram_block1a74.port_b_logical_ram_width = 258;
defparam ram_block1a74.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a74.port_b_read_enable_clock = "clock1";
defparam ram_block1a74.ram_block_type = "auto";

cycloneive_ram_block ram_block1a73(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[73]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a73_PORTBDATAOUT_bus));
defparam ram_block1a73.clk1_output_clock_enable = "ena1";
defparam ram_block1a73.data_interleave_offset_in_bits = 1;
defparam ram_block1a73.data_interleave_width_in_bits = 1;
defparam ram_block1a73.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a73.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a73.operation_mode = "dual_port";
defparam ram_block1a73.port_a_address_clear = "none";
defparam ram_block1a73.port_a_address_width = 3;
defparam ram_block1a73.port_a_data_out_clear = "none";
defparam ram_block1a73.port_a_data_out_clock = "none";
defparam ram_block1a73.port_a_data_width = 1;
defparam ram_block1a73.port_a_first_address = 0;
defparam ram_block1a73.port_a_first_bit_number = 73;
defparam ram_block1a73.port_a_last_address = 7;
defparam ram_block1a73.port_a_logical_ram_depth = 8;
defparam ram_block1a73.port_a_logical_ram_width = 258;
defparam ram_block1a73.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a73.port_b_address_clear = "none";
defparam ram_block1a73.port_b_address_clock = "clock1";
defparam ram_block1a73.port_b_address_width = 3;
defparam ram_block1a73.port_b_data_out_clear = "none";
defparam ram_block1a73.port_b_data_out_clock = "clock1";
defparam ram_block1a73.port_b_data_width = 1;
defparam ram_block1a73.port_b_first_address = 0;
defparam ram_block1a73.port_b_first_bit_number = 73;
defparam ram_block1a73.port_b_last_address = 7;
defparam ram_block1a73.port_b_logical_ram_depth = 8;
defparam ram_block1a73.port_b_logical_ram_width = 258;
defparam ram_block1a73.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a73.port_b_read_enable_clock = "clock1";
defparam ram_block1a73.ram_block_type = "auto";

cycloneive_ram_block ram_block1a72(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[72]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a72_PORTBDATAOUT_bus));
defparam ram_block1a72.clk1_output_clock_enable = "ena1";
defparam ram_block1a72.data_interleave_offset_in_bits = 1;
defparam ram_block1a72.data_interleave_width_in_bits = 1;
defparam ram_block1a72.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a72.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a72.operation_mode = "dual_port";
defparam ram_block1a72.port_a_address_clear = "none";
defparam ram_block1a72.port_a_address_width = 3;
defparam ram_block1a72.port_a_data_out_clear = "none";
defparam ram_block1a72.port_a_data_out_clock = "none";
defparam ram_block1a72.port_a_data_width = 1;
defparam ram_block1a72.port_a_first_address = 0;
defparam ram_block1a72.port_a_first_bit_number = 72;
defparam ram_block1a72.port_a_last_address = 7;
defparam ram_block1a72.port_a_logical_ram_depth = 8;
defparam ram_block1a72.port_a_logical_ram_width = 258;
defparam ram_block1a72.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a72.port_b_address_clear = "none";
defparam ram_block1a72.port_b_address_clock = "clock1";
defparam ram_block1a72.port_b_address_width = 3;
defparam ram_block1a72.port_b_data_out_clear = "none";
defparam ram_block1a72.port_b_data_out_clock = "clock1";
defparam ram_block1a72.port_b_data_width = 1;
defparam ram_block1a72.port_b_first_address = 0;
defparam ram_block1a72.port_b_first_bit_number = 72;
defparam ram_block1a72.port_b_last_address = 7;
defparam ram_block1a72.port_b_logical_ram_depth = 8;
defparam ram_block1a72.port_b_logical_ram_width = 258;
defparam ram_block1a72.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a72.port_b_read_enable_clock = "clock1";
defparam ram_block1a72.ram_block_type = "auto";

cycloneive_ram_block ram_block1a71(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[71]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a71_PORTBDATAOUT_bus));
defparam ram_block1a71.clk1_output_clock_enable = "ena1";
defparam ram_block1a71.data_interleave_offset_in_bits = 1;
defparam ram_block1a71.data_interleave_width_in_bits = 1;
defparam ram_block1a71.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a71.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a71.operation_mode = "dual_port";
defparam ram_block1a71.port_a_address_clear = "none";
defparam ram_block1a71.port_a_address_width = 3;
defparam ram_block1a71.port_a_data_out_clear = "none";
defparam ram_block1a71.port_a_data_out_clock = "none";
defparam ram_block1a71.port_a_data_width = 1;
defparam ram_block1a71.port_a_first_address = 0;
defparam ram_block1a71.port_a_first_bit_number = 71;
defparam ram_block1a71.port_a_last_address = 7;
defparam ram_block1a71.port_a_logical_ram_depth = 8;
defparam ram_block1a71.port_a_logical_ram_width = 258;
defparam ram_block1a71.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a71.port_b_address_clear = "none";
defparam ram_block1a71.port_b_address_clock = "clock1";
defparam ram_block1a71.port_b_address_width = 3;
defparam ram_block1a71.port_b_data_out_clear = "none";
defparam ram_block1a71.port_b_data_out_clock = "clock1";
defparam ram_block1a71.port_b_data_width = 1;
defparam ram_block1a71.port_b_first_address = 0;
defparam ram_block1a71.port_b_first_bit_number = 71;
defparam ram_block1a71.port_b_last_address = 7;
defparam ram_block1a71.port_b_logical_ram_depth = 8;
defparam ram_block1a71.port_b_logical_ram_width = 258;
defparam ram_block1a71.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a71.port_b_read_enable_clock = "clock1";
defparam ram_block1a71.ram_block_type = "auto";

cycloneive_ram_block ram_block1a70(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[70]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a70_PORTBDATAOUT_bus));
defparam ram_block1a70.clk1_output_clock_enable = "ena1";
defparam ram_block1a70.data_interleave_offset_in_bits = 1;
defparam ram_block1a70.data_interleave_width_in_bits = 1;
defparam ram_block1a70.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a70.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a70.operation_mode = "dual_port";
defparam ram_block1a70.port_a_address_clear = "none";
defparam ram_block1a70.port_a_address_width = 3;
defparam ram_block1a70.port_a_data_out_clear = "none";
defparam ram_block1a70.port_a_data_out_clock = "none";
defparam ram_block1a70.port_a_data_width = 1;
defparam ram_block1a70.port_a_first_address = 0;
defparam ram_block1a70.port_a_first_bit_number = 70;
defparam ram_block1a70.port_a_last_address = 7;
defparam ram_block1a70.port_a_logical_ram_depth = 8;
defparam ram_block1a70.port_a_logical_ram_width = 258;
defparam ram_block1a70.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a70.port_b_address_clear = "none";
defparam ram_block1a70.port_b_address_clock = "clock1";
defparam ram_block1a70.port_b_address_width = 3;
defparam ram_block1a70.port_b_data_out_clear = "none";
defparam ram_block1a70.port_b_data_out_clock = "clock1";
defparam ram_block1a70.port_b_data_width = 1;
defparam ram_block1a70.port_b_first_address = 0;
defparam ram_block1a70.port_b_first_bit_number = 70;
defparam ram_block1a70.port_b_last_address = 7;
defparam ram_block1a70.port_b_logical_ram_depth = 8;
defparam ram_block1a70.port_b_logical_ram_width = 258;
defparam ram_block1a70.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a70.port_b_read_enable_clock = "clock1";
defparam ram_block1a70.ram_block_type = "auto";

cycloneive_ram_block ram_block1a69(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[69]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a69_PORTBDATAOUT_bus));
defparam ram_block1a69.clk1_output_clock_enable = "ena1";
defparam ram_block1a69.data_interleave_offset_in_bits = 1;
defparam ram_block1a69.data_interleave_width_in_bits = 1;
defparam ram_block1a69.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a69.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a69.operation_mode = "dual_port";
defparam ram_block1a69.port_a_address_clear = "none";
defparam ram_block1a69.port_a_address_width = 3;
defparam ram_block1a69.port_a_data_out_clear = "none";
defparam ram_block1a69.port_a_data_out_clock = "none";
defparam ram_block1a69.port_a_data_width = 1;
defparam ram_block1a69.port_a_first_address = 0;
defparam ram_block1a69.port_a_first_bit_number = 69;
defparam ram_block1a69.port_a_last_address = 7;
defparam ram_block1a69.port_a_logical_ram_depth = 8;
defparam ram_block1a69.port_a_logical_ram_width = 258;
defparam ram_block1a69.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a69.port_b_address_clear = "none";
defparam ram_block1a69.port_b_address_clock = "clock1";
defparam ram_block1a69.port_b_address_width = 3;
defparam ram_block1a69.port_b_data_out_clear = "none";
defparam ram_block1a69.port_b_data_out_clock = "clock1";
defparam ram_block1a69.port_b_data_width = 1;
defparam ram_block1a69.port_b_first_address = 0;
defparam ram_block1a69.port_b_first_bit_number = 69;
defparam ram_block1a69.port_b_last_address = 7;
defparam ram_block1a69.port_b_logical_ram_depth = 8;
defparam ram_block1a69.port_b_logical_ram_width = 258;
defparam ram_block1a69.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a69.port_b_read_enable_clock = "clock1";
defparam ram_block1a69.ram_block_type = "auto";

cycloneive_ram_block ram_block1a68(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[68]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a68_PORTBDATAOUT_bus));
defparam ram_block1a68.clk1_output_clock_enable = "ena1";
defparam ram_block1a68.data_interleave_offset_in_bits = 1;
defparam ram_block1a68.data_interleave_width_in_bits = 1;
defparam ram_block1a68.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a68.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a68.operation_mode = "dual_port";
defparam ram_block1a68.port_a_address_clear = "none";
defparam ram_block1a68.port_a_address_width = 3;
defparam ram_block1a68.port_a_data_out_clear = "none";
defparam ram_block1a68.port_a_data_out_clock = "none";
defparam ram_block1a68.port_a_data_width = 1;
defparam ram_block1a68.port_a_first_address = 0;
defparam ram_block1a68.port_a_first_bit_number = 68;
defparam ram_block1a68.port_a_last_address = 7;
defparam ram_block1a68.port_a_logical_ram_depth = 8;
defparam ram_block1a68.port_a_logical_ram_width = 258;
defparam ram_block1a68.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a68.port_b_address_clear = "none";
defparam ram_block1a68.port_b_address_clock = "clock1";
defparam ram_block1a68.port_b_address_width = 3;
defparam ram_block1a68.port_b_data_out_clear = "none";
defparam ram_block1a68.port_b_data_out_clock = "clock1";
defparam ram_block1a68.port_b_data_width = 1;
defparam ram_block1a68.port_b_first_address = 0;
defparam ram_block1a68.port_b_first_bit_number = 68;
defparam ram_block1a68.port_b_last_address = 7;
defparam ram_block1a68.port_b_logical_ram_depth = 8;
defparam ram_block1a68.port_b_logical_ram_width = 258;
defparam ram_block1a68.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a68.port_b_read_enable_clock = "clock1";
defparam ram_block1a68.ram_block_type = "auto";

cycloneive_ram_block ram_block1a138(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[138]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a138_PORTBDATAOUT_bus));
defparam ram_block1a138.clk1_output_clock_enable = "ena1";
defparam ram_block1a138.data_interleave_offset_in_bits = 1;
defparam ram_block1a138.data_interleave_width_in_bits = 1;
defparam ram_block1a138.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a138.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a138.operation_mode = "dual_port";
defparam ram_block1a138.port_a_address_clear = "none";
defparam ram_block1a138.port_a_address_width = 3;
defparam ram_block1a138.port_a_data_out_clear = "none";
defparam ram_block1a138.port_a_data_out_clock = "none";
defparam ram_block1a138.port_a_data_width = 1;
defparam ram_block1a138.port_a_first_address = 0;
defparam ram_block1a138.port_a_first_bit_number = 138;
defparam ram_block1a138.port_a_last_address = 7;
defparam ram_block1a138.port_a_logical_ram_depth = 8;
defparam ram_block1a138.port_a_logical_ram_width = 258;
defparam ram_block1a138.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a138.port_b_address_clear = "none";
defparam ram_block1a138.port_b_address_clock = "clock1";
defparam ram_block1a138.port_b_address_width = 3;
defparam ram_block1a138.port_b_data_out_clear = "none";
defparam ram_block1a138.port_b_data_out_clock = "clock1";
defparam ram_block1a138.port_b_data_width = 1;
defparam ram_block1a138.port_b_first_address = 0;
defparam ram_block1a138.port_b_first_bit_number = 138;
defparam ram_block1a138.port_b_last_address = 7;
defparam ram_block1a138.port_b_logical_ram_depth = 8;
defparam ram_block1a138.port_b_logical_ram_width = 258;
defparam ram_block1a138.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a138.port_b_read_enable_clock = "clock1";
defparam ram_block1a138.ram_block_type = "auto";

cycloneive_ram_block ram_block1a137(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[137]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a137_PORTBDATAOUT_bus));
defparam ram_block1a137.clk1_output_clock_enable = "ena1";
defparam ram_block1a137.data_interleave_offset_in_bits = 1;
defparam ram_block1a137.data_interleave_width_in_bits = 1;
defparam ram_block1a137.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a137.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a137.operation_mode = "dual_port";
defparam ram_block1a137.port_a_address_clear = "none";
defparam ram_block1a137.port_a_address_width = 3;
defparam ram_block1a137.port_a_data_out_clear = "none";
defparam ram_block1a137.port_a_data_out_clock = "none";
defparam ram_block1a137.port_a_data_width = 1;
defparam ram_block1a137.port_a_first_address = 0;
defparam ram_block1a137.port_a_first_bit_number = 137;
defparam ram_block1a137.port_a_last_address = 7;
defparam ram_block1a137.port_a_logical_ram_depth = 8;
defparam ram_block1a137.port_a_logical_ram_width = 258;
defparam ram_block1a137.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a137.port_b_address_clear = "none";
defparam ram_block1a137.port_b_address_clock = "clock1";
defparam ram_block1a137.port_b_address_width = 3;
defparam ram_block1a137.port_b_data_out_clear = "none";
defparam ram_block1a137.port_b_data_out_clock = "clock1";
defparam ram_block1a137.port_b_data_width = 1;
defparam ram_block1a137.port_b_first_address = 0;
defparam ram_block1a137.port_b_first_bit_number = 137;
defparam ram_block1a137.port_b_last_address = 7;
defparam ram_block1a137.port_b_logical_ram_depth = 8;
defparam ram_block1a137.port_b_logical_ram_width = 258;
defparam ram_block1a137.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a137.port_b_read_enable_clock = "clock1";
defparam ram_block1a137.ram_block_type = "auto";

cycloneive_ram_block ram_block1a136(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[136]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a136_PORTBDATAOUT_bus));
defparam ram_block1a136.clk1_output_clock_enable = "ena1";
defparam ram_block1a136.data_interleave_offset_in_bits = 1;
defparam ram_block1a136.data_interleave_width_in_bits = 1;
defparam ram_block1a136.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a136.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a136.operation_mode = "dual_port";
defparam ram_block1a136.port_a_address_clear = "none";
defparam ram_block1a136.port_a_address_width = 3;
defparam ram_block1a136.port_a_data_out_clear = "none";
defparam ram_block1a136.port_a_data_out_clock = "none";
defparam ram_block1a136.port_a_data_width = 1;
defparam ram_block1a136.port_a_first_address = 0;
defparam ram_block1a136.port_a_first_bit_number = 136;
defparam ram_block1a136.port_a_last_address = 7;
defparam ram_block1a136.port_a_logical_ram_depth = 8;
defparam ram_block1a136.port_a_logical_ram_width = 258;
defparam ram_block1a136.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a136.port_b_address_clear = "none";
defparam ram_block1a136.port_b_address_clock = "clock1";
defparam ram_block1a136.port_b_address_width = 3;
defparam ram_block1a136.port_b_data_out_clear = "none";
defparam ram_block1a136.port_b_data_out_clock = "clock1";
defparam ram_block1a136.port_b_data_width = 1;
defparam ram_block1a136.port_b_first_address = 0;
defparam ram_block1a136.port_b_first_bit_number = 136;
defparam ram_block1a136.port_b_last_address = 7;
defparam ram_block1a136.port_b_logical_ram_depth = 8;
defparam ram_block1a136.port_b_logical_ram_width = 258;
defparam ram_block1a136.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a136.port_b_read_enable_clock = "clock1";
defparam ram_block1a136.ram_block_type = "auto";

cycloneive_ram_block ram_block1a135(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[135]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a135_PORTBDATAOUT_bus));
defparam ram_block1a135.clk1_output_clock_enable = "ena1";
defparam ram_block1a135.data_interleave_offset_in_bits = 1;
defparam ram_block1a135.data_interleave_width_in_bits = 1;
defparam ram_block1a135.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a135.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a135.operation_mode = "dual_port";
defparam ram_block1a135.port_a_address_clear = "none";
defparam ram_block1a135.port_a_address_width = 3;
defparam ram_block1a135.port_a_data_out_clear = "none";
defparam ram_block1a135.port_a_data_out_clock = "none";
defparam ram_block1a135.port_a_data_width = 1;
defparam ram_block1a135.port_a_first_address = 0;
defparam ram_block1a135.port_a_first_bit_number = 135;
defparam ram_block1a135.port_a_last_address = 7;
defparam ram_block1a135.port_a_logical_ram_depth = 8;
defparam ram_block1a135.port_a_logical_ram_width = 258;
defparam ram_block1a135.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a135.port_b_address_clear = "none";
defparam ram_block1a135.port_b_address_clock = "clock1";
defparam ram_block1a135.port_b_address_width = 3;
defparam ram_block1a135.port_b_data_out_clear = "none";
defparam ram_block1a135.port_b_data_out_clock = "clock1";
defparam ram_block1a135.port_b_data_width = 1;
defparam ram_block1a135.port_b_first_address = 0;
defparam ram_block1a135.port_b_first_bit_number = 135;
defparam ram_block1a135.port_b_last_address = 7;
defparam ram_block1a135.port_b_logical_ram_depth = 8;
defparam ram_block1a135.port_b_logical_ram_width = 258;
defparam ram_block1a135.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a135.port_b_read_enable_clock = "clock1";
defparam ram_block1a135.ram_block_type = "auto";

cycloneive_ram_block ram_block1a134(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[134]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a134_PORTBDATAOUT_bus));
defparam ram_block1a134.clk1_output_clock_enable = "ena1";
defparam ram_block1a134.data_interleave_offset_in_bits = 1;
defparam ram_block1a134.data_interleave_width_in_bits = 1;
defparam ram_block1a134.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a134.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a134.operation_mode = "dual_port";
defparam ram_block1a134.port_a_address_clear = "none";
defparam ram_block1a134.port_a_address_width = 3;
defparam ram_block1a134.port_a_data_out_clear = "none";
defparam ram_block1a134.port_a_data_out_clock = "none";
defparam ram_block1a134.port_a_data_width = 1;
defparam ram_block1a134.port_a_first_address = 0;
defparam ram_block1a134.port_a_first_bit_number = 134;
defparam ram_block1a134.port_a_last_address = 7;
defparam ram_block1a134.port_a_logical_ram_depth = 8;
defparam ram_block1a134.port_a_logical_ram_width = 258;
defparam ram_block1a134.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a134.port_b_address_clear = "none";
defparam ram_block1a134.port_b_address_clock = "clock1";
defparam ram_block1a134.port_b_address_width = 3;
defparam ram_block1a134.port_b_data_out_clear = "none";
defparam ram_block1a134.port_b_data_out_clock = "clock1";
defparam ram_block1a134.port_b_data_width = 1;
defparam ram_block1a134.port_b_first_address = 0;
defparam ram_block1a134.port_b_first_bit_number = 134;
defparam ram_block1a134.port_b_last_address = 7;
defparam ram_block1a134.port_b_logical_ram_depth = 8;
defparam ram_block1a134.port_b_logical_ram_width = 258;
defparam ram_block1a134.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a134.port_b_read_enable_clock = "clock1";
defparam ram_block1a134.ram_block_type = "auto";

cycloneive_ram_block ram_block1a133(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[133]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a133_PORTBDATAOUT_bus));
defparam ram_block1a133.clk1_output_clock_enable = "ena1";
defparam ram_block1a133.data_interleave_offset_in_bits = 1;
defparam ram_block1a133.data_interleave_width_in_bits = 1;
defparam ram_block1a133.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a133.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a133.operation_mode = "dual_port";
defparam ram_block1a133.port_a_address_clear = "none";
defparam ram_block1a133.port_a_address_width = 3;
defparam ram_block1a133.port_a_data_out_clear = "none";
defparam ram_block1a133.port_a_data_out_clock = "none";
defparam ram_block1a133.port_a_data_width = 1;
defparam ram_block1a133.port_a_first_address = 0;
defparam ram_block1a133.port_a_first_bit_number = 133;
defparam ram_block1a133.port_a_last_address = 7;
defparam ram_block1a133.port_a_logical_ram_depth = 8;
defparam ram_block1a133.port_a_logical_ram_width = 258;
defparam ram_block1a133.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a133.port_b_address_clear = "none";
defparam ram_block1a133.port_b_address_clock = "clock1";
defparam ram_block1a133.port_b_address_width = 3;
defparam ram_block1a133.port_b_data_out_clear = "none";
defparam ram_block1a133.port_b_data_out_clock = "clock1";
defparam ram_block1a133.port_b_data_width = 1;
defparam ram_block1a133.port_b_first_address = 0;
defparam ram_block1a133.port_b_first_bit_number = 133;
defparam ram_block1a133.port_b_last_address = 7;
defparam ram_block1a133.port_b_logical_ram_depth = 8;
defparam ram_block1a133.port_b_logical_ram_width = 258;
defparam ram_block1a133.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a133.port_b_read_enable_clock = "clock1";
defparam ram_block1a133.ram_block_type = "auto";

cycloneive_ram_block ram_block1a132(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[132]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a132_PORTBDATAOUT_bus));
defparam ram_block1a132.clk1_output_clock_enable = "ena1";
defparam ram_block1a132.data_interleave_offset_in_bits = 1;
defparam ram_block1a132.data_interleave_width_in_bits = 1;
defparam ram_block1a132.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a132.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a132.operation_mode = "dual_port";
defparam ram_block1a132.port_a_address_clear = "none";
defparam ram_block1a132.port_a_address_width = 3;
defparam ram_block1a132.port_a_data_out_clear = "none";
defparam ram_block1a132.port_a_data_out_clock = "none";
defparam ram_block1a132.port_a_data_width = 1;
defparam ram_block1a132.port_a_first_address = 0;
defparam ram_block1a132.port_a_first_bit_number = 132;
defparam ram_block1a132.port_a_last_address = 7;
defparam ram_block1a132.port_a_logical_ram_depth = 8;
defparam ram_block1a132.port_a_logical_ram_width = 258;
defparam ram_block1a132.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a132.port_b_address_clear = "none";
defparam ram_block1a132.port_b_address_clock = "clock1";
defparam ram_block1a132.port_b_address_width = 3;
defparam ram_block1a132.port_b_data_out_clear = "none";
defparam ram_block1a132.port_b_data_out_clock = "clock1";
defparam ram_block1a132.port_b_data_width = 1;
defparam ram_block1a132.port_b_first_address = 0;
defparam ram_block1a132.port_b_first_bit_number = 132;
defparam ram_block1a132.port_b_last_address = 7;
defparam ram_block1a132.port_b_logical_ram_depth = 8;
defparam ram_block1a132.port_b_logical_ram_width = 258;
defparam ram_block1a132.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a132.port_b_read_enable_clock = "clock1";
defparam ram_block1a132.ram_block_type = "auto";

cycloneive_ram_block ram_block1a202(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[202]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a202_PORTBDATAOUT_bus));
defparam ram_block1a202.clk1_output_clock_enable = "ena1";
defparam ram_block1a202.data_interleave_offset_in_bits = 1;
defparam ram_block1a202.data_interleave_width_in_bits = 1;
defparam ram_block1a202.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a202.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a202.operation_mode = "dual_port";
defparam ram_block1a202.port_a_address_clear = "none";
defparam ram_block1a202.port_a_address_width = 3;
defparam ram_block1a202.port_a_data_out_clear = "none";
defparam ram_block1a202.port_a_data_out_clock = "none";
defparam ram_block1a202.port_a_data_width = 1;
defparam ram_block1a202.port_a_first_address = 0;
defparam ram_block1a202.port_a_first_bit_number = 202;
defparam ram_block1a202.port_a_last_address = 7;
defparam ram_block1a202.port_a_logical_ram_depth = 8;
defparam ram_block1a202.port_a_logical_ram_width = 258;
defparam ram_block1a202.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a202.port_b_address_clear = "none";
defparam ram_block1a202.port_b_address_clock = "clock1";
defparam ram_block1a202.port_b_address_width = 3;
defparam ram_block1a202.port_b_data_out_clear = "none";
defparam ram_block1a202.port_b_data_out_clock = "clock1";
defparam ram_block1a202.port_b_data_width = 1;
defparam ram_block1a202.port_b_first_address = 0;
defparam ram_block1a202.port_b_first_bit_number = 202;
defparam ram_block1a202.port_b_last_address = 7;
defparam ram_block1a202.port_b_logical_ram_depth = 8;
defparam ram_block1a202.port_b_logical_ram_width = 258;
defparam ram_block1a202.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a202.port_b_read_enable_clock = "clock1";
defparam ram_block1a202.ram_block_type = "auto";

cycloneive_ram_block ram_block1a201(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[201]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a201_PORTBDATAOUT_bus));
defparam ram_block1a201.clk1_output_clock_enable = "ena1";
defparam ram_block1a201.data_interleave_offset_in_bits = 1;
defparam ram_block1a201.data_interleave_width_in_bits = 1;
defparam ram_block1a201.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a201.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a201.operation_mode = "dual_port";
defparam ram_block1a201.port_a_address_clear = "none";
defparam ram_block1a201.port_a_address_width = 3;
defparam ram_block1a201.port_a_data_out_clear = "none";
defparam ram_block1a201.port_a_data_out_clock = "none";
defparam ram_block1a201.port_a_data_width = 1;
defparam ram_block1a201.port_a_first_address = 0;
defparam ram_block1a201.port_a_first_bit_number = 201;
defparam ram_block1a201.port_a_last_address = 7;
defparam ram_block1a201.port_a_logical_ram_depth = 8;
defparam ram_block1a201.port_a_logical_ram_width = 258;
defparam ram_block1a201.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a201.port_b_address_clear = "none";
defparam ram_block1a201.port_b_address_clock = "clock1";
defparam ram_block1a201.port_b_address_width = 3;
defparam ram_block1a201.port_b_data_out_clear = "none";
defparam ram_block1a201.port_b_data_out_clock = "clock1";
defparam ram_block1a201.port_b_data_width = 1;
defparam ram_block1a201.port_b_first_address = 0;
defparam ram_block1a201.port_b_first_bit_number = 201;
defparam ram_block1a201.port_b_last_address = 7;
defparam ram_block1a201.port_b_logical_ram_depth = 8;
defparam ram_block1a201.port_b_logical_ram_width = 258;
defparam ram_block1a201.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a201.port_b_read_enable_clock = "clock1";
defparam ram_block1a201.ram_block_type = "auto";

cycloneive_ram_block ram_block1a200(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[200]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a200_PORTBDATAOUT_bus));
defparam ram_block1a200.clk1_output_clock_enable = "ena1";
defparam ram_block1a200.data_interleave_offset_in_bits = 1;
defparam ram_block1a200.data_interleave_width_in_bits = 1;
defparam ram_block1a200.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a200.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a200.operation_mode = "dual_port";
defparam ram_block1a200.port_a_address_clear = "none";
defparam ram_block1a200.port_a_address_width = 3;
defparam ram_block1a200.port_a_data_out_clear = "none";
defparam ram_block1a200.port_a_data_out_clock = "none";
defparam ram_block1a200.port_a_data_width = 1;
defparam ram_block1a200.port_a_first_address = 0;
defparam ram_block1a200.port_a_first_bit_number = 200;
defparam ram_block1a200.port_a_last_address = 7;
defparam ram_block1a200.port_a_logical_ram_depth = 8;
defparam ram_block1a200.port_a_logical_ram_width = 258;
defparam ram_block1a200.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a200.port_b_address_clear = "none";
defparam ram_block1a200.port_b_address_clock = "clock1";
defparam ram_block1a200.port_b_address_width = 3;
defparam ram_block1a200.port_b_data_out_clear = "none";
defparam ram_block1a200.port_b_data_out_clock = "clock1";
defparam ram_block1a200.port_b_data_width = 1;
defparam ram_block1a200.port_b_first_address = 0;
defparam ram_block1a200.port_b_first_bit_number = 200;
defparam ram_block1a200.port_b_last_address = 7;
defparam ram_block1a200.port_b_logical_ram_depth = 8;
defparam ram_block1a200.port_b_logical_ram_width = 258;
defparam ram_block1a200.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a200.port_b_read_enable_clock = "clock1";
defparam ram_block1a200.ram_block_type = "auto";

cycloneive_ram_block ram_block1a199(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[199]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a199_PORTBDATAOUT_bus));
defparam ram_block1a199.clk1_output_clock_enable = "ena1";
defparam ram_block1a199.data_interleave_offset_in_bits = 1;
defparam ram_block1a199.data_interleave_width_in_bits = 1;
defparam ram_block1a199.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a199.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a199.operation_mode = "dual_port";
defparam ram_block1a199.port_a_address_clear = "none";
defparam ram_block1a199.port_a_address_width = 3;
defparam ram_block1a199.port_a_data_out_clear = "none";
defparam ram_block1a199.port_a_data_out_clock = "none";
defparam ram_block1a199.port_a_data_width = 1;
defparam ram_block1a199.port_a_first_address = 0;
defparam ram_block1a199.port_a_first_bit_number = 199;
defparam ram_block1a199.port_a_last_address = 7;
defparam ram_block1a199.port_a_logical_ram_depth = 8;
defparam ram_block1a199.port_a_logical_ram_width = 258;
defparam ram_block1a199.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a199.port_b_address_clear = "none";
defparam ram_block1a199.port_b_address_clock = "clock1";
defparam ram_block1a199.port_b_address_width = 3;
defparam ram_block1a199.port_b_data_out_clear = "none";
defparam ram_block1a199.port_b_data_out_clock = "clock1";
defparam ram_block1a199.port_b_data_width = 1;
defparam ram_block1a199.port_b_first_address = 0;
defparam ram_block1a199.port_b_first_bit_number = 199;
defparam ram_block1a199.port_b_last_address = 7;
defparam ram_block1a199.port_b_logical_ram_depth = 8;
defparam ram_block1a199.port_b_logical_ram_width = 258;
defparam ram_block1a199.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a199.port_b_read_enable_clock = "clock1";
defparam ram_block1a199.ram_block_type = "auto";

cycloneive_ram_block ram_block1a198(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[198]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a198_PORTBDATAOUT_bus));
defparam ram_block1a198.clk1_output_clock_enable = "ena1";
defparam ram_block1a198.data_interleave_offset_in_bits = 1;
defparam ram_block1a198.data_interleave_width_in_bits = 1;
defparam ram_block1a198.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a198.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a198.operation_mode = "dual_port";
defparam ram_block1a198.port_a_address_clear = "none";
defparam ram_block1a198.port_a_address_width = 3;
defparam ram_block1a198.port_a_data_out_clear = "none";
defparam ram_block1a198.port_a_data_out_clock = "none";
defparam ram_block1a198.port_a_data_width = 1;
defparam ram_block1a198.port_a_first_address = 0;
defparam ram_block1a198.port_a_first_bit_number = 198;
defparam ram_block1a198.port_a_last_address = 7;
defparam ram_block1a198.port_a_logical_ram_depth = 8;
defparam ram_block1a198.port_a_logical_ram_width = 258;
defparam ram_block1a198.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a198.port_b_address_clear = "none";
defparam ram_block1a198.port_b_address_clock = "clock1";
defparam ram_block1a198.port_b_address_width = 3;
defparam ram_block1a198.port_b_data_out_clear = "none";
defparam ram_block1a198.port_b_data_out_clock = "clock1";
defparam ram_block1a198.port_b_data_width = 1;
defparam ram_block1a198.port_b_first_address = 0;
defparam ram_block1a198.port_b_first_bit_number = 198;
defparam ram_block1a198.port_b_last_address = 7;
defparam ram_block1a198.port_b_logical_ram_depth = 8;
defparam ram_block1a198.port_b_logical_ram_width = 258;
defparam ram_block1a198.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a198.port_b_read_enable_clock = "clock1";
defparam ram_block1a198.ram_block_type = "auto";

cycloneive_ram_block ram_block1a197(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[197]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a197_PORTBDATAOUT_bus));
defparam ram_block1a197.clk1_output_clock_enable = "ena1";
defparam ram_block1a197.data_interleave_offset_in_bits = 1;
defparam ram_block1a197.data_interleave_width_in_bits = 1;
defparam ram_block1a197.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a197.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a197.operation_mode = "dual_port";
defparam ram_block1a197.port_a_address_clear = "none";
defparam ram_block1a197.port_a_address_width = 3;
defparam ram_block1a197.port_a_data_out_clear = "none";
defparam ram_block1a197.port_a_data_out_clock = "none";
defparam ram_block1a197.port_a_data_width = 1;
defparam ram_block1a197.port_a_first_address = 0;
defparam ram_block1a197.port_a_first_bit_number = 197;
defparam ram_block1a197.port_a_last_address = 7;
defparam ram_block1a197.port_a_logical_ram_depth = 8;
defparam ram_block1a197.port_a_logical_ram_width = 258;
defparam ram_block1a197.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a197.port_b_address_clear = "none";
defparam ram_block1a197.port_b_address_clock = "clock1";
defparam ram_block1a197.port_b_address_width = 3;
defparam ram_block1a197.port_b_data_out_clear = "none";
defparam ram_block1a197.port_b_data_out_clock = "clock1";
defparam ram_block1a197.port_b_data_width = 1;
defparam ram_block1a197.port_b_first_address = 0;
defparam ram_block1a197.port_b_first_bit_number = 197;
defparam ram_block1a197.port_b_last_address = 7;
defparam ram_block1a197.port_b_logical_ram_depth = 8;
defparam ram_block1a197.port_b_logical_ram_width = 258;
defparam ram_block1a197.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a197.port_b_read_enable_clock = "clock1";
defparam ram_block1a197.ram_block_type = "auto";

cycloneive_ram_block ram_block1a196(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[196]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a196_PORTBDATAOUT_bus));
defparam ram_block1a196.clk1_output_clock_enable = "ena1";
defparam ram_block1a196.data_interleave_offset_in_bits = 1;
defparam ram_block1a196.data_interleave_width_in_bits = 1;
defparam ram_block1a196.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a196.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a196.operation_mode = "dual_port";
defparam ram_block1a196.port_a_address_clear = "none";
defparam ram_block1a196.port_a_address_width = 3;
defparam ram_block1a196.port_a_data_out_clear = "none";
defparam ram_block1a196.port_a_data_out_clock = "none";
defparam ram_block1a196.port_a_data_width = 1;
defparam ram_block1a196.port_a_first_address = 0;
defparam ram_block1a196.port_a_first_bit_number = 196;
defparam ram_block1a196.port_a_last_address = 7;
defparam ram_block1a196.port_a_logical_ram_depth = 8;
defparam ram_block1a196.port_a_logical_ram_width = 258;
defparam ram_block1a196.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a196.port_b_address_clear = "none";
defparam ram_block1a196.port_b_address_clock = "clock1";
defparam ram_block1a196.port_b_address_width = 3;
defparam ram_block1a196.port_b_data_out_clear = "none";
defparam ram_block1a196.port_b_data_out_clock = "clock1";
defparam ram_block1a196.port_b_data_width = 1;
defparam ram_block1a196.port_b_first_address = 0;
defparam ram_block1a196.port_b_first_bit_number = 196;
defparam ram_block1a196.port_b_last_address = 7;
defparam ram_block1a196.port_b_logical_ram_depth = 8;
defparam ram_block1a196.port_b_logical_ram_width = 258;
defparam ram_block1a196.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a196.port_b_read_enable_clock = "clock1";
defparam ram_block1a196.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 258;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 258;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 258;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 258;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 258;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 258;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 258;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 258;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 258;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 258;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 258;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 258;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 258;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 258;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a107(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[107]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a107_PORTBDATAOUT_bus));
defparam ram_block1a107.clk1_output_clock_enable = "ena1";
defparam ram_block1a107.data_interleave_offset_in_bits = 1;
defparam ram_block1a107.data_interleave_width_in_bits = 1;
defparam ram_block1a107.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a107.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a107.operation_mode = "dual_port";
defparam ram_block1a107.port_a_address_clear = "none";
defparam ram_block1a107.port_a_address_width = 3;
defparam ram_block1a107.port_a_data_out_clear = "none";
defparam ram_block1a107.port_a_data_out_clock = "none";
defparam ram_block1a107.port_a_data_width = 1;
defparam ram_block1a107.port_a_first_address = 0;
defparam ram_block1a107.port_a_first_bit_number = 107;
defparam ram_block1a107.port_a_last_address = 7;
defparam ram_block1a107.port_a_logical_ram_depth = 8;
defparam ram_block1a107.port_a_logical_ram_width = 258;
defparam ram_block1a107.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a107.port_b_address_clear = "none";
defparam ram_block1a107.port_b_address_clock = "clock1";
defparam ram_block1a107.port_b_address_width = 3;
defparam ram_block1a107.port_b_data_out_clear = "none";
defparam ram_block1a107.port_b_data_out_clock = "clock1";
defparam ram_block1a107.port_b_data_width = 1;
defparam ram_block1a107.port_b_first_address = 0;
defparam ram_block1a107.port_b_first_bit_number = 107;
defparam ram_block1a107.port_b_last_address = 7;
defparam ram_block1a107.port_b_logical_ram_depth = 8;
defparam ram_block1a107.port_b_logical_ram_width = 258;
defparam ram_block1a107.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a107.port_b_read_enable_clock = "clock1";
defparam ram_block1a107.ram_block_type = "auto";

cycloneive_ram_block ram_block1a123(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[123]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a123_PORTBDATAOUT_bus));
defparam ram_block1a123.clk1_output_clock_enable = "ena1";
defparam ram_block1a123.data_interleave_offset_in_bits = 1;
defparam ram_block1a123.data_interleave_width_in_bits = 1;
defparam ram_block1a123.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a123.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a123.operation_mode = "dual_port";
defparam ram_block1a123.port_a_address_clear = "none";
defparam ram_block1a123.port_a_address_width = 3;
defparam ram_block1a123.port_a_data_out_clear = "none";
defparam ram_block1a123.port_a_data_out_clock = "none";
defparam ram_block1a123.port_a_data_width = 1;
defparam ram_block1a123.port_a_first_address = 0;
defparam ram_block1a123.port_a_first_bit_number = 123;
defparam ram_block1a123.port_a_last_address = 7;
defparam ram_block1a123.port_a_logical_ram_depth = 8;
defparam ram_block1a123.port_a_logical_ram_width = 258;
defparam ram_block1a123.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a123.port_b_address_clear = "none";
defparam ram_block1a123.port_b_address_clock = "clock1";
defparam ram_block1a123.port_b_address_width = 3;
defparam ram_block1a123.port_b_data_out_clear = "none";
defparam ram_block1a123.port_b_data_out_clock = "clock1";
defparam ram_block1a123.port_b_data_width = 1;
defparam ram_block1a123.port_b_first_address = 0;
defparam ram_block1a123.port_b_first_bit_number = 123;
defparam ram_block1a123.port_b_last_address = 7;
defparam ram_block1a123.port_b_logical_ram_depth = 8;
defparam ram_block1a123.port_b_logical_ram_width = 258;
defparam ram_block1a123.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a123.port_b_read_enable_clock = "clock1";
defparam ram_block1a123.ram_block_type = "auto";

cycloneive_ram_block ram_block1a91(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[91]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a91_PORTBDATAOUT_bus));
defparam ram_block1a91.clk1_output_clock_enable = "ena1";
defparam ram_block1a91.data_interleave_offset_in_bits = 1;
defparam ram_block1a91.data_interleave_width_in_bits = 1;
defparam ram_block1a91.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a91.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a91.operation_mode = "dual_port";
defparam ram_block1a91.port_a_address_clear = "none";
defparam ram_block1a91.port_a_address_width = 3;
defparam ram_block1a91.port_a_data_out_clear = "none";
defparam ram_block1a91.port_a_data_out_clock = "none";
defparam ram_block1a91.port_a_data_width = 1;
defparam ram_block1a91.port_a_first_address = 0;
defparam ram_block1a91.port_a_first_bit_number = 91;
defparam ram_block1a91.port_a_last_address = 7;
defparam ram_block1a91.port_a_logical_ram_depth = 8;
defparam ram_block1a91.port_a_logical_ram_width = 258;
defparam ram_block1a91.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a91.port_b_address_clear = "none";
defparam ram_block1a91.port_b_address_clock = "clock1";
defparam ram_block1a91.port_b_address_width = 3;
defparam ram_block1a91.port_b_data_out_clear = "none";
defparam ram_block1a91.port_b_data_out_clock = "clock1";
defparam ram_block1a91.port_b_data_width = 1;
defparam ram_block1a91.port_b_first_address = 0;
defparam ram_block1a91.port_b_first_bit_number = 91;
defparam ram_block1a91.port_b_last_address = 7;
defparam ram_block1a91.port_b_logical_ram_depth = 8;
defparam ram_block1a91.port_b_logical_ram_width = 258;
defparam ram_block1a91.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a91.port_b_read_enable_clock = "clock1";
defparam ram_block1a91.ram_block_type = "auto";

cycloneive_ram_block ram_block1a75(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[75]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a75_PORTBDATAOUT_bus));
defparam ram_block1a75.clk1_output_clock_enable = "ena1";
defparam ram_block1a75.data_interleave_offset_in_bits = 1;
defparam ram_block1a75.data_interleave_width_in_bits = 1;
defparam ram_block1a75.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a75.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a75.operation_mode = "dual_port";
defparam ram_block1a75.port_a_address_clear = "none";
defparam ram_block1a75.port_a_address_width = 3;
defparam ram_block1a75.port_a_data_out_clear = "none";
defparam ram_block1a75.port_a_data_out_clock = "none";
defparam ram_block1a75.port_a_data_width = 1;
defparam ram_block1a75.port_a_first_address = 0;
defparam ram_block1a75.port_a_first_bit_number = 75;
defparam ram_block1a75.port_a_last_address = 7;
defparam ram_block1a75.port_a_logical_ram_depth = 8;
defparam ram_block1a75.port_a_logical_ram_width = 258;
defparam ram_block1a75.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a75.port_b_address_clear = "none";
defparam ram_block1a75.port_b_address_clock = "clock1";
defparam ram_block1a75.port_b_address_width = 3;
defparam ram_block1a75.port_b_data_out_clear = "none";
defparam ram_block1a75.port_b_data_out_clock = "clock1";
defparam ram_block1a75.port_b_data_width = 1;
defparam ram_block1a75.port_b_first_address = 0;
defparam ram_block1a75.port_b_first_bit_number = 75;
defparam ram_block1a75.port_b_last_address = 7;
defparam ram_block1a75.port_b_logical_ram_depth = 8;
defparam ram_block1a75.port_b_logical_ram_width = 258;
defparam ram_block1a75.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a75.port_b_read_enable_clock = "clock1";
defparam ram_block1a75.ram_block_type = "auto";

cycloneive_ram_block ram_block1a171(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[171]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a171_PORTBDATAOUT_bus));
defparam ram_block1a171.clk1_output_clock_enable = "ena1";
defparam ram_block1a171.data_interleave_offset_in_bits = 1;
defparam ram_block1a171.data_interleave_width_in_bits = 1;
defparam ram_block1a171.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a171.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a171.operation_mode = "dual_port";
defparam ram_block1a171.port_a_address_clear = "none";
defparam ram_block1a171.port_a_address_width = 3;
defparam ram_block1a171.port_a_data_out_clear = "none";
defparam ram_block1a171.port_a_data_out_clock = "none";
defparam ram_block1a171.port_a_data_width = 1;
defparam ram_block1a171.port_a_first_address = 0;
defparam ram_block1a171.port_a_first_bit_number = 171;
defparam ram_block1a171.port_a_last_address = 7;
defparam ram_block1a171.port_a_logical_ram_depth = 8;
defparam ram_block1a171.port_a_logical_ram_width = 258;
defparam ram_block1a171.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a171.port_b_address_clear = "none";
defparam ram_block1a171.port_b_address_clock = "clock1";
defparam ram_block1a171.port_b_address_width = 3;
defparam ram_block1a171.port_b_data_out_clear = "none";
defparam ram_block1a171.port_b_data_out_clock = "clock1";
defparam ram_block1a171.port_b_data_width = 1;
defparam ram_block1a171.port_b_first_address = 0;
defparam ram_block1a171.port_b_first_bit_number = 171;
defparam ram_block1a171.port_b_last_address = 7;
defparam ram_block1a171.port_b_logical_ram_depth = 8;
defparam ram_block1a171.port_b_logical_ram_width = 258;
defparam ram_block1a171.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a171.port_b_read_enable_clock = "clock1";
defparam ram_block1a171.ram_block_type = "auto";

cycloneive_ram_block ram_block1a187(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[187]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a187_PORTBDATAOUT_bus));
defparam ram_block1a187.clk1_output_clock_enable = "ena1";
defparam ram_block1a187.data_interleave_offset_in_bits = 1;
defparam ram_block1a187.data_interleave_width_in_bits = 1;
defparam ram_block1a187.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a187.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a187.operation_mode = "dual_port";
defparam ram_block1a187.port_a_address_clear = "none";
defparam ram_block1a187.port_a_address_width = 3;
defparam ram_block1a187.port_a_data_out_clear = "none";
defparam ram_block1a187.port_a_data_out_clock = "none";
defparam ram_block1a187.port_a_data_width = 1;
defparam ram_block1a187.port_a_first_address = 0;
defparam ram_block1a187.port_a_first_bit_number = 187;
defparam ram_block1a187.port_a_last_address = 7;
defparam ram_block1a187.port_a_logical_ram_depth = 8;
defparam ram_block1a187.port_a_logical_ram_width = 258;
defparam ram_block1a187.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a187.port_b_address_clear = "none";
defparam ram_block1a187.port_b_address_clock = "clock1";
defparam ram_block1a187.port_b_address_width = 3;
defparam ram_block1a187.port_b_data_out_clear = "none";
defparam ram_block1a187.port_b_data_out_clock = "clock1";
defparam ram_block1a187.port_b_data_width = 1;
defparam ram_block1a187.port_b_first_address = 0;
defparam ram_block1a187.port_b_first_bit_number = 187;
defparam ram_block1a187.port_b_last_address = 7;
defparam ram_block1a187.port_b_logical_ram_depth = 8;
defparam ram_block1a187.port_b_logical_ram_width = 258;
defparam ram_block1a187.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a187.port_b_read_enable_clock = "clock1";
defparam ram_block1a187.ram_block_type = "auto";

cycloneive_ram_block ram_block1a155(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[155]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a155_PORTBDATAOUT_bus));
defparam ram_block1a155.clk1_output_clock_enable = "ena1";
defparam ram_block1a155.data_interleave_offset_in_bits = 1;
defparam ram_block1a155.data_interleave_width_in_bits = 1;
defparam ram_block1a155.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a155.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a155.operation_mode = "dual_port";
defparam ram_block1a155.port_a_address_clear = "none";
defparam ram_block1a155.port_a_address_width = 3;
defparam ram_block1a155.port_a_data_out_clear = "none";
defparam ram_block1a155.port_a_data_out_clock = "none";
defparam ram_block1a155.port_a_data_width = 1;
defparam ram_block1a155.port_a_first_address = 0;
defparam ram_block1a155.port_a_first_bit_number = 155;
defparam ram_block1a155.port_a_last_address = 7;
defparam ram_block1a155.port_a_logical_ram_depth = 8;
defparam ram_block1a155.port_a_logical_ram_width = 258;
defparam ram_block1a155.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a155.port_b_address_clear = "none";
defparam ram_block1a155.port_b_address_clock = "clock1";
defparam ram_block1a155.port_b_address_width = 3;
defparam ram_block1a155.port_b_data_out_clear = "none";
defparam ram_block1a155.port_b_data_out_clock = "clock1";
defparam ram_block1a155.port_b_data_width = 1;
defparam ram_block1a155.port_b_first_address = 0;
defparam ram_block1a155.port_b_first_bit_number = 155;
defparam ram_block1a155.port_b_last_address = 7;
defparam ram_block1a155.port_b_logical_ram_depth = 8;
defparam ram_block1a155.port_b_logical_ram_width = 258;
defparam ram_block1a155.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a155.port_b_read_enable_clock = "clock1";
defparam ram_block1a155.ram_block_type = "auto";

cycloneive_ram_block ram_block1a139(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[139]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a139_PORTBDATAOUT_bus));
defparam ram_block1a139.clk1_output_clock_enable = "ena1";
defparam ram_block1a139.data_interleave_offset_in_bits = 1;
defparam ram_block1a139.data_interleave_width_in_bits = 1;
defparam ram_block1a139.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a139.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a139.operation_mode = "dual_port";
defparam ram_block1a139.port_a_address_clear = "none";
defparam ram_block1a139.port_a_address_width = 3;
defparam ram_block1a139.port_a_data_out_clear = "none";
defparam ram_block1a139.port_a_data_out_clock = "none";
defparam ram_block1a139.port_a_data_width = 1;
defparam ram_block1a139.port_a_first_address = 0;
defparam ram_block1a139.port_a_first_bit_number = 139;
defparam ram_block1a139.port_a_last_address = 7;
defparam ram_block1a139.port_a_logical_ram_depth = 8;
defparam ram_block1a139.port_a_logical_ram_width = 258;
defparam ram_block1a139.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a139.port_b_address_clear = "none";
defparam ram_block1a139.port_b_address_clock = "clock1";
defparam ram_block1a139.port_b_address_width = 3;
defparam ram_block1a139.port_b_data_out_clear = "none";
defparam ram_block1a139.port_b_data_out_clock = "clock1";
defparam ram_block1a139.port_b_data_width = 1;
defparam ram_block1a139.port_b_first_address = 0;
defparam ram_block1a139.port_b_first_bit_number = 139;
defparam ram_block1a139.port_b_last_address = 7;
defparam ram_block1a139.port_b_logical_ram_depth = 8;
defparam ram_block1a139.port_b_logical_ram_width = 258;
defparam ram_block1a139.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a139.port_b_read_enable_clock = "clock1";
defparam ram_block1a139.ram_block_type = "auto";

cycloneive_ram_block ram_block1a235(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[235]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a235_PORTBDATAOUT_bus));
defparam ram_block1a235.clk1_output_clock_enable = "ena1";
defparam ram_block1a235.data_interleave_offset_in_bits = 1;
defparam ram_block1a235.data_interleave_width_in_bits = 1;
defparam ram_block1a235.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a235.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a235.operation_mode = "dual_port";
defparam ram_block1a235.port_a_address_clear = "none";
defparam ram_block1a235.port_a_address_width = 3;
defparam ram_block1a235.port_a_data_out_clear = "none";
defparam ram_block1a235.port_a_data_out_clock = "none";
defparam ram_block1a235.port_a_data_width = 1;
defparam ram_block1a235.port_a_first_address = 0;
defparam ram_block1a235.port_a_first_bit_number = 235;
defparam ram_block1a235.port_a_last_address = 7;
defparam ram_block1a235.port_a_logical_ram_depth = 8;
defparam ram_block1a235.port_a_logical_ram_width = 258;
defparam ram_block1a235.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a235.port_b_address_clear = "none";
defparam ram_block1a235.port_b_address_clock = "clock1";
defparam ram_block1a235.port_b_address_width = 3;
defparam ram_block1a235.port_b_data_out_clear = "none";
defparam ram_block1a235.port_b_data_out_clock = "clock1";
defparam ram_block1a235.port_b_data_width = 1;
defparam ram_block1a235.port_b_first_address = 0;
defparam ram_block1a235.port_b_first_bit_number = 235;
defparam ram_block1a235.port_b_last_address = 7;
defparam ram_block1a235.port_b_logical_ram_depth = 8;
defparam ram_block1a235.port_b_logical_ram_width = 258;
defparam ram_block1a235.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a235.port_b_read_enable_clock = "clock1";
defparam ram_block1a235.ram_block_type = "auto";

cycloneive_ram_block ram_block1a251(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[251]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a251_PORTBDATAOUT_bus));
defparam ram_block1a251.clk1_output_clock_enable = "ena1";
defparam ram_block1a251.data_interleave_offset_in_bits = 1;
defparam ram_block1a251.data_interleave_width_in_bits = 1;
defparam ram_block1a251.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a251.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a251.operation_mode = "dual_port";
defparam ram_block1a251.port_a_address_clear = "none";
defparam ram_block1a251.port_a_address_width = 3;
defparam ram_block1a251.port_a_data_out_clear = "none";
defparam ram_block1a251.port_a_data_out_clock = "none";
defparam ram_block1a251.port_a_data_width = 1;
defparam ram_block1a251.port_a_first_address = 0;
defparam ram_block1a251.port_a_first_bit_number = 251;
defparam ram_block1a251.port_a_last_address = 7;
defparam ram_block1a251.port_a_logical_ram_depth = 8;
defparam ram_block1a251.port_a_logical_ram_width = 258;
defparam ram_block1a251.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a251.port_b_address_clear = "none";
defparam ram_block1a251.port_b_address_clock = "clock1";
defparam ram_block1a251.port_b_address_width = 3;
defparam ram_block1a251.port_b_data_out_clear = "none";
defparam ram_block1a251.port_b_data_out_clock = "clock1";
defparam ram_block1a251.port_b_data_width = 1;
defparam ram_block1a251.port_b_first_address = 0;
defparam ram_block1a251.port_b_first_bit_number = 251;
defparam ram_block1a251.port_b_last_address = 7;
defparam ram_block1a251.port_b_logical_ram_depth = 8;
defparam ram_block1a251.port_b_logical_ram_width = 258;
defparam ram_block1a251.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a251.port_b_read_enable_clock = "clock1";
defparam ram_block1a251.ram_block_type = "auto";

cycloneive_ram_block ram_block1a219(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[219]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a219_PORTBDATAOUT_bus));
defparam ram_block1a219.clk1_output_clock_enable = "ena1";
defparam ram_block1a219.data_interleave_offset_in_bits = 1;
defparam ram_block1a219.data_interleave_width_in_bits = 1;
defparam ram_block1a219.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a219.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a219.operation_mode = "dual_port";
defparam ram_block1a219.port_a_address_clear = "none";
defparam ram_block1a219.port_a_address_width = 3;
defparam ram_block1a219.port_a_data_out_clear = "none";
defparam ram_block1a219.port_a_data_out_clock = "none";
defparam ram_block1a219.port_a_data_width = 1;
defparam ram_block1a219.port_a_first_address = 0;
defparam ram_block1a219.port_a_first_bit_number = 219;
defparam ram_block1a219.port_a_last_address = 7;
defparam ram_block1a219.port_a_logical_ram_depth = 8;
defparam ram_block1a219.port_a_logical_ram_width = 258;
defparam ram_block1a219.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a219.port_b_address_clear = "none";
defparam ram_block1a219.port_b_address_clock = "clock1";
defparam ram_block1a219.port_b_address_width = 3;
defparam ram_block1a219.port_b_data_out_clear = "none";
defparam ram_block1a219.port_b_data_out_clock = "clock1";
defparam ram_block1a219.port_b_data_width = 1;
defparam ram_block1a219.port_b_first_address = 0;
defparam ram_block1a219.port_b_first_bit_number = 219;
defparam ram_block1a219.port_b_last_address = 7;
defparam ram_block1a219.port_b_logical_ram_depth = 8;
defparam ram_block1a219.port_b_logical_ram_width = 258;
defparam ram_block1a219.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a219.port_b_read_enable_clock = "clock1";
defparam ram_block1a219.ram_block_type = "auto";

cycloneive_ram_block ram_block1a203(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[203]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a203_PORTBDATAOUT_bus));
defparam ram_block1a203.clk1_output_clock_enable = "ena1";
defparam ram_block1a203.data_interleave_offset_in_bits = 1;
defparam ram_block1a203.data_interleave_width_in_bits = 1;
defparam ram_block1a203.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a203.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a203.operation_mode = "dual_port";
defparam ram_block1a203.port_a_address_clear = "none";
defparam ram_block1a203.port_a_address_width = 3;
defparam ram_block1a203.port_a_data_out_clear = "none";
defparam ram_block1a203.port_a_data_out_clock = "none";
defparam ram_block1a203.port_a_data_width = 1;
defparam ram_block1a203.port_a_first_address = 0;
defparam ram_block1a203.port_a_first_bit_number = 203;
defparam ram_block1a203.port_a_last_address = 7;
defparam ram_block1a203.port_a_logical_ram_depth = 8;
defparam ram_block1a203.port_a_logical_ram_width = 258;
defparam ram_block1a203.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a203.port_b_address_clear = "none";
defparam ram_block1a203.port_b_address_clock = "clock1";
defparam ram_block1a203.port_b_address_width = 3;
defparam ram_block1a203.port_b_data_out_clear = "none";
defparam ram_block1a203.port_b_data_out_clock = "clock1";
defparam ram_block1a203.port_b_data_width = 1;
defparam ram_block1a203.port_b_first_address = 0;
defparam ram_block1a203.port_b_first_bit_number = 203;
defparam ram_block1a203.port_b_last_address = 7;
defparam ram_block1a203.port_b_logical_ram_depth = 8;
defparam ram_block1a203.port_b_logical_ram_width = 258;
defparam ram_block1a203.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a203.port_b_read_enable_clock = "clock1";
defparam ram_block1a203.ram_block_type = "auto";

cycloneive_ram_block ram_block1a43(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[43]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a43_PORTBDATAOUT_bus));
defparam ram_block1a43.clk1_output_clock_enable = "ena1";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a43.operation_mode = "dual_port";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 3;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "none";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 0;
defparam ram_block1a43.port_a_first_bit_number = 43;
defparam ram_block1a43.port_a_last_address = 7;
defparam ram_block1a43.port_a_logical_ram_depth = 8;
defparam ram_block1a43.port_a_logical_ram_width = 258;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a43.port_b_address_clear = "none";
defparam ram_block1a43.port_b_address_clock = "clock1";
defparam ram_block1a43.port_b_address_width = 3;
defparam ram_block1a43.port_b_data_out_clear = "none";
defparam ram_block1a43.port_b_data_out_clock = "clock1";
defparam ram_block1a43.port_b_data_width = 1;
defparam ram_block1a43.port_b_first_address = 0;
defparam ram_block1a43.port_b_first_bit_number = 43;
defparam ram_block1a43.port_b_last_address = 7;
defparam ram_block1a43.port_b_logical_ram_depth = 8;
defparam ram_block1a43.port_b_logical_ram_width = 258;
defparam ram_block1a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a43.port_b_read_enable_clock = "clock1";
defparam ram_block1a43.ram_block_type = "auto";

cycloneive_ram_block ram_block1a59(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[59]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a59_PORTBDATAOUT_bus));
defparam ram_block1a59.clk1_output_clock_enable = "ena1";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a59.operation_mode = "dual_port";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 3;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "none";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 0;
defparam ram_block1a59.port_a_first_bit_number = 59;
defparam ram_block1a59.port_a_last_address = 7;
defparam ram_block1a59.port_a_logical_ram_depth = 8;
defparam ram_block1a59.port_a_logical_ram_width = 258;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a59.port_b_address_clear = "none";
defparam ram_block1a59.port_b_address_clock = "clock1";
defparam ram_block1a59.port_b_address_width = 3;
defparam ram_block1a59.port_b_data_out_clear = "none";
defparam ram_block1a59.port_b_data_out_clock = "clock1";
defparam ram_block1a59.port_b_data_width = 1;
defparam ram_block1a59.port_b_first_address = 0;
defparam ram_block1a59.port_b_first_bit_number = 59;
defparam ram_block1a59.port_b_last_address = 7;
defparam ram_block1a59.port_b_logical_ram_depth = 8;
defparam ram_block1a59.port_b_logical_ram_width = 258;
defparam ram_block1a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a59.port_b_read_enable_clock = "clock1";
defparam ram_block1a59.ram_block_type = "auto";

cycloneive_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk1_output_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 3;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 7;
defparam ram_block1a27.port_a_logical_ram_depth = 8;
defparam ram_block1a27.port_a_logical_ram_width = 258;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 3;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock1";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 7;
defparam ram_block1a27.port_b_logical_ram_depth = 8;
defparam ram_block1a27.port_b_logical_ram_width = 258;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 258;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 258;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a108(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[108]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a108_PORTBDATAOUT_bus));
defparam ram_block1a108.clk1_output_clock_enable = "ena1";
defparam ram_block1a108.data_interleave_offset_in_bits = 1;
defparam ram_block1a108.data_interleave_width_in_bits = 1;
defparam ram_block1a108.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a108.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a108.operation_mode = "dual_port";
defparam ram_block1a108.port_a_address_clear = "none";
defparam ram_block1a108.port_a_address_width = 3;
defparam ram_block1a108.port_a_data_out_clear = "none";
defparam ram_block1a108.port_a_data_out_clock = "none";
defparam ram_block1a108.port_a_data_width = 1;
defparam ram_block1a108.port_a_first_address = 0;
defparam ram_block1a108.port_a_first_bit_number = 108;
defparam ram_block1a108.port_a_last_address = 7;
defparam ram_block1a108.port_a_logical_ram_depth = 8;
defparam ram_block1a108.port_a_logical_ram_width = 258;
defparam ram_block1a108.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a108.port_b_address_clear = "none";
defparam ram_block1a108.port_b_address_clock = "clock1";
defparam ram_block1a108.port_b_address_width = 3;
defparam ram_block1a108.port_b_data_out_clear = "none";
defparam ram_block1a108.port_b_data_out_clock = "clock1";
defparam ram_block1a108.port_b_data_width = 1;
defparam ram_block1a108.port_b_first_address = 0;
defparam ram_block1a108.port_b_first_bit_number = 108;
defparam ram_block1a108.port_b_last_address = 7;
defparam ram_block1a108.port_b_logical_ram_depth = 8;
defparam ram_block1a108.port_b_logical_ram_width = 258;
defparam ram_block1a108.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a108.port_b_read_enable_clock = "clock1";
defparam ram_block1a108.ram_block_type = "auto";

cycloneive_ram_block ram_block1a172(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[172]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a172_PORTBDATAOUT_bus));
defparam ram_block1a172.clk1_output_clock_enable = "ena1";
defparam ram_block1a172.data_interleave_offset_in_bits = 1;
defparam ram_block1a172.data_interleave_width_in_bits = 1;
defparam ram_block1a172.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a172.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a172.operation_mode = "dual_port";
defparam ram_block1a172.port_a_address_clear = "none";
defparam ram_block1a172.port_a_address_width = 3;
defparam ram_block1a172.port_a_data_out_clear = "none";
defparam ram_block1a172.port_a_data_out_clock = "none";
defparam ram_block1a172.port_a_data_width = 1;
defparam ram_block1a172.port_a_first_address = 0;
defparam ram_block1a172.port_a_first_bit_number = 172;
defparam ram_block1a172.port_a_last_address = 7;
defparam ram_block1a172.port_a_logical_ram_depth = 8;
defparam ram_block1a172.port_a_logical_ram_width = 258;
defparam ram_block1a172.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a172.port_b_address_clear = "none";
defparam ram_block1a172.port_b_address_clock = "clock1";
defparam ram_block1a172.port_b_address_width = 3;
defparam ram_block1a172.port_b_data_out_clear = "none";
defparam ram_block1a172.port_b_data_out_clock = "clock1";
defparam ram_block1a172.port_b_data_width = 1;
defparam ram_block1a172.port_b_first_address = 0;
defparam ram_block1a172.port_b_first_bit_number = 172;
defparam ram_block1a172.port_b_last_address = 7;
defparam ram_block1a172.port_b_logical_ram_depth = 8;
defparam ram_block1a172.port_b_logical_ram_width = 258;
defparam ram_block1a172.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a172.port_b_read_enable_clock = "clock1";
defparam ram_block1a172.ram_block_type = "auto";

cycloneive_ram_block ram_block1a236(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[236]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a236_PORTBDATAOUT_bus));
defparam ram_block1a236.clk1_output_clock_enable = "ena1";
defparam ram_block1a236.data_interleave_offset_in_bits = 1;
defparam ram_block1a236.data_interleave_width_in_bits = 1;
defparam ram_block1a236.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a236.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a236.operation_mode = "dual_port";
defparam ram_block1a236.port_a_address_clear = "none";
defparam ram_block1a236.port_a_address_width = 3;
defparam ram_block1a236.port_a_data_out_clear = "none";
defparam ram_block1a236.port_a_data_out_clock = "none";
defparam ram_block1a236.port_a_data_width = 1;
defparam ram_block1a236.port_a_first_address = 0;
defparam ram_block1a236.port_a_first_bit_number = 236;
defparam ram_block1a236.port_a_last_address = 7;
defparam ram_block1a236.port_a_logical_ram_depth = 8;
defparam ram_block1a236.port_a_logical_ram_width = 258;
defparam ram_block1a236.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a236.port_b_address_clear = "none";
defparam ram_block1a236.port_b_address_clock = "clock1";
defparam ram_block1a236.port_b_address_width = 3;
defparam ram_block1a236.port_b_data_out_clear = "none";
defparam ram_block1a236.port_b_data_out_clock = "clock1";
defparam ram_block1a236.port_b_data_width = 1;
defparam ram_block1a236.port_b_first_address = 0;
defparam ram_block1a236.port_b_first_bit_number = 236;
defparam ram_block1a236.port_b_last_address = 7;
defparam ram_block1a236.port_b_logical_ram_depth = 8;
defparam ram_block1a236.port_b_logical_ram_width = 258;
defparam ram_block1a236.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a236.port_b_read_enable_clock = "clock1";
defparam ram_block1a236.ram_block_type = "auto";

cycloneive_ram_block ram_block1a44(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[44]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a44_PORTBDATAOUT_bus));
defparam ram_block1a44.clk1_output_clock_enable = "ena1";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a44.operation_mode = "dual_port";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 3;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "none";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 0;
defparam ram_block1a44.port_a_first_bit_number = 44;
defparam ram_block1a44.port_a_last_address = 7;
defparam ram_block1a44.port_a_logical_ram_depth = 8;
defparam ram_block1a44.port_a_logical_ram_width = 258;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a44.port_b_address_clear = "none";
defparam ram_block1a44.port_b_address_clock = "clock1";
defparam ram_block1a44.port_b_address_width = 3;
defparam ram_block1a44.port_b_data_out_clear = "none";
defparam ram_block1a44.port_b_data_out_clock = "clock1";
defparam ram_block1a44.port_b_data_width = 1;
defparam ram_block1a44.port_b_first_address = 0;
defparam ram_block1a44.port_b_first_bit_number = 44;
defparam ram_block1a44.port_b_last_address = 7;
defparam ram_block1a44.port_b_logical_ram_depth = 8;
defparam ram_block1a44.port_b_logical_ram_width = 258;
defparam ram_block1a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a44.port_b_read_enable_clock = "clock1";
defparam ram_block1a44.ram_block_type = "auto";

cycloneive_ram_block ram_block1a124(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[124]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a124_PORTBDATAOUT_bus));
defparam ram_block1a124.clk1_output_clock_enable = "ena1";
defparam ram_block1a124.data_interleave_offset_in_bits = 1;
defparam ram_block1a124.data_interleave_width_in_bits = 1;
defparam ram_block1a124.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a124.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a124.operation_mode = "dual_port";
defparam ram_block1a124.port_a_address_clear = "none";
defparam ram_block1a124.port_a_address_width = 3;
defparam ram_block1a124.port_a_data_out_clear = "none";
defparam ram_block1a124.port_a_data_out_clock = "none";
defparam ram_block1a124.port_a_data_width = 1;
defparam ram_block1a124.port_a_first_address = 0;
defparam ram_block1a124.port_a_first_bit_number = 124;
defparam ram_block1a124.port_a_last_address = 7;
defparam ram_block1a124.port_a_logical_ram_depth = 8;
defparam ram_block1a124.port_a_logical_ram_width = 258;
defparam ram_block1a124.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a124.port_b_address_clear = "none";
defparam ram_block1a124.port_b_address_clock = "clock1";
defparam ram_block1a124.port_b_address_width = 3;
defparam ram_block1a124.port_b_data_out_clear = "none";
defparam ram_block1a124.port_b_data_out_clock = "clock1";
defparam ram_block1a124.port_b_data_width = 1;
defparam ram_block1a124.port_b_first_address = 0;
defparam ram_block1a124.port_b_first_bit_number = 124;
defparam ram_block1a124.port_b_last_address = 7;
defparam ram_block1a124.port_b_logical_ram_depth = 8;
defparam ram_block1a124.port_b_logical_ram_width = 258;
defparam ram_block1a124.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a124.port_b_read_enable_clock = "clock1";
defparam ram_block1a124.ram_block_type = "auto";

cycloneive_ram_block ram_block1a188(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[188]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a188_PORTBDATAOUT_bus));
defparam ram_block1a188.clk1_output_clock_enable = "ena1";
defparam ram_block1a188.data_interleave_offset_in_bits = 1;
defparam ram_block1a188.data_interleave_width_in_bits = 1;
defparam ram_block1a188.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a188.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a188.operation_mode = "dual_port";
defparam ram_block1a188.port_a_address_clear = "none";
defparam ram_block1a188.port_a_address_width = 3;
defparam ram_block1a188.port_a_data_out_clear = "none";
defparam ram_block1a188.port_a_data_out_clock = "none";
defparam ram_block1a188.port_a_data_width = 1;
defparam ram_block1a188.port_a_first_address = 0;
defparam ram_block1a188.port_a_first_bit_number = 188;
defparam ram_block1a188.port_a_last_address = 7;
defparam ram_block1a188.port_a_logical_ram_depth = 8;
defparam ram_block1a188.port_a_logical_ram_width = 258;
defparam ram_block1a188.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a188.port_b_address_clear = "none";
defparam ram_block1a188.port_b_address_clock = "clock1";
defparam ram_block1a188.port_b_address_width = 3;
defparam ram_block1a188.port_b_data_out_clear = "none";
defparam ram_block1a188.port_b_data_out_clock = "clock1";
defparam ram_block1a188.port_b_data_width = 1;
defparam ram_block1a188.port_b_first_address = 0;
defparam ram_block1a188.port_b_first_bit_number = 188;
defparam ram_block1a188.port_b_last_address = 7;
defparam ram_block1a188.port_b_logical_ram_depth = 8;
defparam ram_block1a188.port_b_logical_ram_width = 258;
defparam ram_block1a188.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a188.port_b_read_enable_clock = "clock1";
defparam ram_block1a188.ram_block_type = "auto";

cycloneive_ram_block ram_block1a252(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[252]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a252_PORTBDATAOUT_bus));
defparam ram_block1a252.clk1_output_clock_enable = "ena1";
defparam ram_block1a252.data_interleave_offset_in_bits = 1;
defparam ram_block1a252.data_interleave_width_in_bits = 1;
defparam ram_block1a252.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a252.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a252.operation_mode = "dual_port";
defparam ram_block1a252.port_a_address_clear = "none";
defparam ram_block1a252.port_a_address_width = 3;
defparam ram_block1a252.port_a_data_out_clear = "none";
defparam ram_block1a252.port_a_data_out_clock = "none";
defparam ram_block1a252.port_a_data_width = 1;
defparam ram_block1a252.port_a_first_address = 0;
defparam ram_block1a252.port_a_first_bit_number = 252;
defparam ram_block1a252.port_a_last_address = 7;
defparam ram_block1a252.port_a_logical_ram_depth = 8;
defparam ram_block1a252.port_a_logical_ram_width = 258;
defparam ram_block1a252.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a252.port_b_address_clear = "none";
defparam ram_block1a252.port_b_address_clock = "clock1";
defparam ram_block1a252.port_b_address_width = 3;
defparam ram_block1a252.port_b_data_out_clear = "none";
defparam ram_block1a252.port_b_data_out_clock = "clock1";
defparam ram_block1a252.port_b_data_width = 1;
defparam ram_block1a252.port_b_first_address = 0;
defparam ram_block1a252.port_b_first_bit_number = 252;
defparam ram_block1a252.port_b_last_address = 7;
defparam ram_block1a252.port_b_logical_ram_depth = 8;
defparam ram_block1a252.port_b_logical_ram_width = 258;
defparam ram_block1a252.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a252.port_b_read_enable_clock = "clock1";
defparam ram_block1a252.ram_block_type = "auto";

cycloneive_ram_block ram_block1a60(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[60]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a60_PORTBDATAOUT_bus));
defparam ram_block1a60.clk1_output_clock_enable = "ena1";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a60.operation_mode = "dual_port";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 3;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "none";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 0;
defparam ram_block1a60.port_a_first_bit_number = 60;
defparam ram_block1a60.port_a_last_address = 7;
defparam ram_block1a60.port_a_logical_ram_depth = 8;
defparam ram_block1a60.port_a_logical_ram_width = 258;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a60.port_b_address_clear = "none";
defparam ram_block1a60.port_b_address_clock = "clock1";
defparam ram_block1a60.port_b_address_width = 3;
defparam ram_block1a60.port_b_data_out_clear = "none";
defparam ram_block1a60.port_b_data_out_clock = "clock1";
defparam ram_block1a60.port_b_data_width = 1;
defparam ram_block1a60.port_b_first_address = 0;
defparam ram_block1a60.port_b_first_bit_number = 60;
defparam ram_block1a60.port_b_last_address = 7;
defparam ram_block1a60.port_b_logical_ram_depth = 8;
defparam ram_block1a60.port_b_logical_ram_width = 258;
defparam ram_block1a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a60.port_b_read_enable_clock = "clock1";
defparam ram_block1a60.ram_block_type = "auto";

cycloneive_ram_block ram_block1a156(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[156]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a156_PORTBDATAOUT_bus));
defparam ram_block1a156.clk1_output_clock_enable = "ena1";
defparam ram_block1a156.data_interleave_offset_in_bits = 1;
defparam ram_block1a156.data_interleave_width_in_bits = 1;
defparam ram_block1a156.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a156.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a156.operation_mode = "dual_port";
defparam ram_block1a156.port_a_address_clear = "none";
defparam ram_block1a156.port_a_address_width = 3;
defparam ram_block1a156.port_a_data_out_clear = "none";
defparam ram_block1a156.port_a_data_out_clock = "none";
defparam ram_block1a156.port_a_data_width = 1;
defparam ram_block1a156.port_a_first_address = 0;
defparam ram_block1a156.port_a_first_bit_number = 156;
defparam ram_block1a156.port_a_last_address = 7;
defparam ram_block1a156.port_a_logical_ram_depth = 8;
defparam ram_block1a156.port_a_logical_ram_width = 258;
defparam ram_block1a156.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a156.port_b_address_clear = "none";
defparam ram_block1a156.port_b_address_clock = "clock1";
defparam ram_block1a156.port_b_address_width = 3;
defparam ram_block1a156.port_b_data_out_clear = "none";
defparam ram_block1a156.port_b_data_out_clock = "clock1";
defparam ram_block1a156.port_b_data_width = 1;
defparam ram_block1a156.port_b_first_address = 0;
defparam ram_block1a156.port_b_first_bit_number = 156;
defparam ram_block1a156.port_b_last_address = 7;
defparam ram_block1a156.port_b_logical_ram_depth = 8;
defparam ram_block1a156.port_b_logical_ram_width = 258;
defparam ram_block1a156.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a156.port_b_read_enable_clock = "clock1";
defparam ram_block1a156.ram_block_type = "auto";

cycloneive_ram_block ram_block1a92(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[92]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a92_PORTBDATAOUT_bus));
defparam ram_block1a92.clk1_output_clock_enable = "ena1";
defparam ram_block1a92.data_interleave_offset_in_bits = 1;
defparam ram_block1a92.data_interleave_width_in_bits = 1;
defparam ram_block1a92.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a92.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a92.operation_mode = "dual_port";
defparam ram_block1a92.port_a_address_clear = "none";
defparam ram_block1a92.port_a_address_width = 3;
defparam ram_block1a92.port_a_data_out_clear = "none";
defparam ram_block1a92.port_a_data_out_clock = "none";
defparam ram_block1a92.port_a_data_width = 1;
defparam ram_block1a92.port_a_first_address = 0;
defparam ram_block1a92.port_a_first_bit_number = 92;
defparam ram_block1a92.port_a_last_address = 7;
defparam ram_block1a92.port_a_logical_ram_depth = 8;
defparam ram_block1a92.port_a_logical_ram_width = 258;
defparam ram_block1a92.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a92.port_b_address_clear = "none";
defparam ram_block1a92.port_b_address_clock = "clock1";
defparam ram_block1a92.port_b_address_width = 3;
defparam ram_block1a92.port_b_data_out_clear = "none";
defparam ram_block1a92.port_b_data_out_clock = "clock1";
defparam ram_block1a92.port_b_data_width = 1;
defparam ram_block1a92.port_b_first_address = 0;
defparam ram_block1a92.port_b_first_bit_number = 92;
defparam ram_block1a92.port_b_last_address = 7;
defparam ram_block1a92.port_b_logical_ram_depth = 8;
defparam ram_block1a92.port_b_logical_ram_width = 258;
defparam ram_block1a92.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a92.port_b_read_enable_clock = "clock1";
defparam ram_block1a92.ram_block_type = "auto";

cycloneive_ram_block ram_block1a220(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[220]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a220_PORTBDATAOUT_bus));
defparam ram_block1a220.clk1_output_clock_enable = "ena1";
defparam ram_block1a220.data_interleave_offset_in_bits = 1;
defparam ram_block1a220.data_interleave_width_in_bits = 1;
defparam ram_block1a220.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a220.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a220.operation_mode = "dual_port";
defparam ram_block1a220.port_a_address_clear = "none";
defparam ram_block1a220.port_a_address_width = 3;
defparam ram_block1a220.port_a_data_out_clear = "none";
defparam ram_block1a220.port_a_data_out_clock = "none";
defparam ram_block1a220.port_a_data_width = 1;
defparam ram_block1a220.port_a_first_address = 0;
defparam ram_block1a220.port_a_first_bit_number = 220;
defparam ram_block1a220.port_a_last_address = 7;
defparam ram_block1a220.port_a_logical_ram_depth = 8;
defparam ram_block1a220.port_a_logical_ram_width = 258;
defparam ram_block1a220.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a220.port_b_address_clear = "none";
defparam ram_block1a220.port_b_address_clock = "clock1";
defparam ram_block1a220.port_b_address_width = 3;
defparam ram_block1a220.port_b_data_out_clear = "none";
defparam ram_block1a220.port_b_data_out_clock = "clock1";
defparam ram_block1a220.port_b_data_width = 1;
defparam ram_block1a220.port_b_first_address = 0;
defparam ram_block1a220.port_b_first_bit_number = 220;
defparam ram_block1a220.port_b_last_address = 7;
defparam ram_block1a220.port_b_logical_ram_depth = 8;
defparam ram_block1a220.port_b_logical_ram_width = 258;
defparam ram_block1a220.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a220.port_b_read_enable_clock = "clock1";
defparam ram_block1a220.ram_block_type = "auto";

cycloneive_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk1_output_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 3;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 7;
defparam ram_block1a28.port_a_logical_ram_depth = 8;
defparam ram_block1a28.port_a_logical_ram_width = 258;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 3;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "clock1";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 7;
defparam ram_block1a28.port_b_logical_ram_depth = 8;
defparam ram_block1a28.port_b_logical_ram_width = 258;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cycloneive_ram_block ram_block1a140(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[140]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a140_PORTBDATAOUT_bus));
defparam ram_block1a140.clk1_output_clock_enable = "ena1";
defparam ram_block1a140.data_interleave_offset_in_bits = 1;
defparam ram_block1a140.data_interleave_width_in_bits = 1;
defparam ram_block1a140.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a140.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a140.operation_mode = "dual_port";
defparam ram_block1a140.port_a_address_clear = "none";
defparam ram_block1a140.port_a_address_width = 3;
defparam ram_block1a140.port_a_data_out_clear = "none";
defparam ram_block1a140.port_a_data_out_clock = "none";
defparam ram_block1a140.port_a_data_width = 1;
defparam ram_block1a140.port_a_first_address = 0;
defparam ram_block1a140.port_a_first_bit_number = 140;
defparam ram_block1a140.port_a_last_address = 7;
defparam ram_block1a140.port_a_logical_ram_depth = 8;
defparam ram_block1a140.port_a_logical_ram_width = 258;
defparam ram_block1a140.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a140.port_b_address_clear = "none";
defparam ram_block1a140.port_b_address_clock = "clock1";
defparam ram_block1a140.port_b_address_width = 3;
defparam ram_block1a140.port_b_data_out_clear = "none";
defparam ram_block1a140.port_b_data_out_clock = "clock1";
defparam ram_block1a140.port_b_data_width = 1;
defparam ram_block1a140.port_b_first_address = 0;
defparam ram_block1a140.port_b_first_bit_number = 140;
defparam ram_block1a140.port_b_last_address = 7;
defparam ram_block1a140.port_b_logical_ram_depth = 8;
defparam ram_block1a140.port_b_logical_ram_width = 258;
defparam ram_block1a140.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a140.port_b_read_enable_clock = "clock1";
defparam ram_block1a140.ram_block_type = "auto";

cycloneive_ram_block ram_block1a76(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[76]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a76_PORTBDATAOUT_bus));
defparam ram_block1a76.clk1_output_clock_enable = "ena1";
defparam ram_block1a76.data_interleave_offset_in_bits = 1;
defparam ram_block1a76.data_interleave_width_in_bits = 1;
defparam ram_block1a76.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a76.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a76.operation_mode = "dual_port";
defparam ram_block1a76.port_a_address_clear = "none";
defparam ram_block1a76.port_a_address_width = 3;
defparam ram_block1a76.port_a_data_out_clear = "none";
defparam ram_block1a76.port_a_data_out_clock = "none";
defparam ram_block1a76.port_a_data_width = 1;
defparam ram_block1a76.port_a_first_address = 0;
defparam ram_block1a76.port_a_first_bit_number = 76;
defparam ram_block1a76.port_a_last_address = 7;
defparam ram_block1a76.port_a_logical_ram_depth = 8;
defparam ram_block1a76.port_a_logical_ram_width = 258;
defparam ram_block1a76.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a76.port_b_address_clear = "none";
defparam ram_block1a76.port_b_address_clock = "clock1";
defparam ram_block1a76.port_b_address_width = 3;
defparam ram_block1a76.port_b_data_out_clear = "none";
defparam ram_block1a76.port_b_data_out_clock = "clock1";
defparam ram_block1a76.port_b_data_width = 1;
defparam ram_block1a76.port_b_first_address = 0;
defparam ram_block1a76.port_b_first_bit_number = 76;
defparam ram_block1a76.port_b_last_address = 7;
defparam ram_block1a76.port_b_logical_ram_depth = 8;
defparam ram_block1a76.port_b_logical_ram_width = 258;
defparam ram_block1a76.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a76.port_b_read_enable_clock = "clock1";
defparam ram_block1a76.ram_block_type = "auto";

cycloneive_ram_block ram_block1a204(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[204]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a204_PORTBDATAOUT_bus));
defparam ram_block1a204.clk1_output_clock_enable = "ena1";
defparam ram_block1a204.data_interleave_offset_in_bits = 1;
defparam ram_block1a204.data_interleave_width_in_bits = 1;
defparam ram_block1a204.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a204.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a204.operation_mode = "dual_port";
defparam ram_block1a204.port_a_address_clear = "none";
defparam ram_block1a204.port_a_address_width = 3;
defparam ram_block1a204.port_a_data_out_clear = "none";
defparam ram_block1a204.port_a_data_out_clock = "none";
defparam ram_block1a204.port_a_data_width = 1;
defparam ram_block1a204.port_a_first_address = 0;
defparam ram_block1a204.port_a_first_bit_number = 204;
defparam ram_block1a204.port_a_last_address = 7;
defparam ram_block1a204.port_a_logical_ram_depth = 8;
defparam ram_block1a204.port_a_logical_ram_width = 258;
defparam ram_block1a204.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a204.port_b_address_clear = "none";
defparam ram_block1a204.port_b_address_clock = "clock1";
defparam ram_block1a204.port_b_address_width = 3;
defparam ram_block1a204.port_b_data_out_clear = "none";
defparam ram_block1a204.port_b_data_out_clock = "clock1";
defparam ram_block1a204.port_b_data_width = 1;
defparam ram_block1a204.port_b_first_address = 0;
defparam ram_block1a204.port_b_first_bit_number = 204;
defparam ram_block1a204.port_b_last_address = 7;
defparam ram_block1a204.port_b_logical_ram_depth = 8;
defparam ram_block1a204.port_b_logical_ram_width = 258;
defparam ram_block1a204.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a204.port_b_read_enable_clock = "clock1";
defparam ram_block1a204.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 258;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 258;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a173(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[173]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a173_PORTBDATAOUT_bus));
defparam ram_block1a173.clk1_output_clock_enable = "ena1";
defparam ram_block1a173.data_interleave_offset_in_bits = 1;
defparam ram_block1a173.data_interleave_width_in_bits = 1;
defparam ram_block1a173.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a173.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a173.operation_mode = "dual_port";
defparam ram_block1a173.port_a_address_clear = "none";
defparam ram_block1a173.port_a_address_width = 3;
defparam ram_block1a173.port_a_data_out_clear = "none";
defparam ram_block1a173.port_a_data_out_clock = "none";
defparam ram_block1a173.port_a_data_width = 1;
defparam ram_block1a173.port_a_first_address = 0;
defparam ram_block1a173.port_a_first_bit_number = 173;
defparam ram_block1a173.port_a_last_address = 7;
defparam ram_block1a173.port_a_logical_ram_depth = 8;
defparam ram_block1a173.port_a_logical_ram_width = 258;
defparam ram_block1a173.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a173.port_b_address_clear = "none";
defparam ram_block1a173.port_b_address_clock = "clock1";
defparam ram_block1a173.port_b_address_width = 3;
defparam ram_block1a173.port_b_data_out_clear = "none";
defparam ram_block1a173.port_b_data_out_clock = "clock1";
defparam ram_block1a173.port_b_data_width = 1;
defparam ram_block1a173.port_b_first_address = 0;
defparam ram_block1a173.port_b_first_bit_number = 173;
defparam ram_block1a173.port_b_last_address = 7;
defparam ram_block1a173.port_b_logical_ram_depth = 8;
defparam ram_block1a173.port_b_logical_ram_width = 258;
defparam ram_block1a173.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a173.port_b_read_enable_clock = "clock1";
defparam ram_block1a173.ram_block_type = "auto";

cycloneive_ram_block ram_block1a189(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[189]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a189_PORTBDATAOUT_bus));
defparam ram_block1a189.clk1_output_clock_enable = "ena1";
defparam ram_block1a189.data_interleave_offset_in_bits = 1;
defparam ram_block1a189.data_interleave_width_in_bits = 1;
defparam ram_block1a189.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a189.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a189.operation_mode = "dual_port";
defparam ram_block1a189.port_a_address_clear = "none";
defparam ram_block1a189.port_a_address_width = 3;
defparam ram_block1a189.port_a_data_out_clear = "none";
defparam ram_block1a189.port_a_data_out_clock = "none";
defparam ram_block1a189.port_a_data_width = 1;
defparam ram_block1a189.port_a_first_address = 0;
defparam ram_block1a189.port_a_first_bit_number = 189;
defparam ram_block1a189.port_a_last_address = 7;
defparam ram_block1a189.port_a_logical_ram_depth = 8;
defparam ram_block1a189.port_a_logical_ram_width = 258;
defparam ram_block1a189.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a189.port_b_address_clear = "none";
defparam ram_block1a189.port_b_address_clock = "clock1";
defparam ram_block1a189.port_b_address_width = 3;
defparam ram_block1a189.port_b_data_out_clear = "none";
defparam ram_block1a189.port_b_data_out_clock = "clock1";
defparam ram_block1a189.port_b_data_width = 1;
defparam ram_block1a189.port_b_first_address = 0;
defparam ram_block1a189.port_b_first_bit_number = 189;
defparam ram_block1a189.port_b_last_address = 7;
defparam ram_block1a189.port_b_logical_ram_depth = 8;
defparam ram_block1a189.port_b_logical_ram_width = 258;
defparam ram_block1a189.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a189.port_b_read_enable_clock = "clock1";
defparam ram_block1a189.ram_block_type = "auto";

cycloneive_ram_block ram_block1a157(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[157]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a157_PORTBDATAOUT_bus));
defparam ram_block1a157.clk1_output_clock_enable = "ena1";
defparam ram_block1a157.data_interleave_offset_in_bits = 1;
defparam ram_block1a157.data_interleave_width_in_bits = 1;
defparam ram_block1a157.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a157.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a157.operation_mode = "dual_port";
defparam ram_block1a157.port_a_address_clear = "none";
defparam ram_block1a157.port_a_address_width = 3;
defparam ram_block1a157.port_a_data_out_clear = "none";
defparam ram_block1a157.port_a_data_out_clock = "none";
defparam ram_block1a157.port_a_data_width = 1;
defparam ram_block1a157.port_a_first_address = 0;
defparam ram_block1a157.port_a_first_bit_number = 157;
defparam ram_block1a157.port_a_last_address = 7;
defparam ram_block1a157.port_a_logical_ram_depth = 8;
defparam ram_block1a157.port_a_logical_ram_width = 258;
defparam ram_block1a157.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a157.port_b_address_clear = "none";
defparam ram_block1a157.port_b_address_clock = "clock1";
defparam ram_block1a157.port_b_address_width = 3;
defparam ram_block1a157.port_b_data_out_clear = "none";
defparam ram_block1a157.port_b_data_out_clock = "clock1";
defparam ram_block1a157.port_b_data_width = 1;
defparam ram_block1a157.port_b_first_address = 0;
defparam ram_block1a157.port_b_first_bit_number = 157;
defparam ram_block1a157.port_b_last_address = 7;
defparam ram_block1a157.port_b_logical_ram_depth = 8;
defparam ram_block1a157.port_b_logical_ram_width = 258;
defparam ram_block1a157.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a157.port_b_read_enable_clock = "clock1";
defparam ram_block1a157.ram_block_type = "auto";

cycloneive_ram_block ram_block1a141(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[141]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a141_PORTBDATAOUT_bus));
defparam ram_block1a141.clk1_output_clock_enable = "ena1";
defparam ram_block1a141.data_interleave_offset_in_bits = 1;
defparam ram_block1a141.data_interleave_width_in_bits = 1;
defparam ram_block1a141.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a141.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a141.operation_mode = "dual_port";
defparam ram_block1a141.port_a_address_clear = "none";
defparam ram_block1a141.port_a_address_width = 3;
defparam ram_block1a141.port_a_data_out_clear = "none";
defparam ram_block1a141.port_a_data_out_clock = "none";
defparam ram_block1a141.port_a_data_width = 1;
defparam ram_block1a141.port_a_first_address = 0;
defparam ram_block1a141.port_a_first_bit_number = 141;
defparam ram_block1a141.port_a_last_address = 7;
defparam ram_block1a141.port_a_logical_ram_depth = 8;
defparam ram_block1a141.port_a_logical_ram_width = 258;
defparam ram_block1a141.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a141.port_b_address_clear = "none";
defparam ram_block1a141.port_b_address_clock = "clock1";
defparam ram_block1a141.port_b_address_width = 3;
defparam ram_block1a141.port_b_data_out_clear = "none";
defparam ram_block1a141.port_b_data_out_clock = "clock1";
defparam ram_block1a141.port_b_data_width = 1;
defparam ram_block1a141.port_b_first_address = 0;
defparam ram_block1a141.port_b_first_bit_number = 141;
defparam ram_block1a141.port_b_last_address = 7;
defparam ram_block1a141.port_b_logical_ram_depth = 8;
defparam ram_block1a141.port_b_logical_ram_width = 258;
defparam ram_block1a141.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a141.port_b_read_enable_clock = "clock1";
defparam ram_block1a141.ram_block_type = "auto";

cycloneive_ram_block ram_block1a109(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[109]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a109_PORTBDATAOUT_bus));
defparam ram_block1a109.clk1_output_clock_enable = "ena1";
defparam ram_block1a109.data_interleave_offset_in_bits = 1;
defparam ram_block1a109.data_interleave_width_in_bits = 1;
defparam ram_block1a109.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a109.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a109.operation_mode = "dual_port";
defparam ram_block1a109.port_a_address_clear = "none";
defparam ram_block1a109.port_a_address_width = 3;
defparam ram_block1a109.port_a_data_out_clear = "none";
defparam ram_block1a109.port_a_data_out_clock = "none";
defparam ram_block1a109.port_a_data_width = 1;
defparam ram_block1a109.port_a_first_address = 0;
defparam ram_block1a109.port_a_first_bit_number = 109;
defparam ram_block1a109.port_a_last_address = 7;
defparam ram_block1a109.port_a_logical_ram_depth = 8;
defparam ram_block1a109.port_a_logical_ram_width = 258;
defparam ram_block1a109.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a109.port_b_address_clear = "none";
defparam ram_block1a109.port_b_address_clock = "clock1";
defparam ram_block1a109.port_b_address_width = 3;
defparam ram_block1a109.port_b_data_out_clear = "none";
defparam ram_block1a109.port_b_data_out_clock = "clock1";
defparam ram_block1a109.port_b_data_width = 1;
defparam ram_block1a109.port_b_first_address = 0;
defparam ram_block1a109.port_b_first_bit_number = 109;
defparam ram_block1a109.port_b_last_address = 7;
defparam ram_block1a109.port_b_logical_ram_depth = 8;
defparam ram_block1a109.port_b_logical_ram_width = 258;
defparam ram_block1a109.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a109.port_b_read_enable_clock = "clock1";
defparam ram_block1a109.ram_block_type = "auto";

cycloneive_ram_block ram_block1a125(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[125]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a125_PORTBDATAOUT_bus));
defparam ram_block1a125.clk1_output_clock_enable = "ena1";
defparam ram_block1a125.data_interleave_offset_in_bits = 1;
defparam ram_block1a125.data_interleave_width_in_bits = 1;
defparam ram_block1a125.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a125.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a125.operation_mode = "dual_port";
defparam ram_block1a125.port_a_address_clear = "none";
defparam ram_block1a125.port_a_address_width = 3;
defparam ram_block1a125.port_a_data_out_clear = "none";
defparam ram_block1a125.port_a_data_out_clock = "none";
defparam ram_block1a125.port_a_data_width = 1;
defparam ram_block1a125.port_a_first_address = 0;
defparam ram_block1a125.port_a_first_bit_number = 125;
defparam ram_block1a125.port_a_last_address = 7;
defparam ram_block1a125.port_a_logical_ram_depth = 8;
defparam ram_block1a125.port_a_logical_ram_width = 258;
defparam ram_block1a125.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a125.port_b_address_clear = "none";
defparam ram_block1a125.port_b_address_clock = "clock1";
defparam ram_block1a125.port_b_address_width = 3;
defparam ram_block1a125.port_b_data_out_clear = "none";
defparam ram_block1a125.port_b_data_out_clock = "clock1";
defparam ram_block1a125.port_b_data_width = 1;
defparam ram_block1a125.port_b_first_address = 0;
defparam ram_block1a125.port_b_first_bit_number = 125;
defparam ram_block1a125.port_b_last_address = 7;
defparam ram_block1a125.port_b_logical_ram_depth = 8;
defparam ram_block1a125.port_b_logical_ram_width = 258;
defparam ram_block1a125.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a125.port_b_read_enable_clock = "clock1";
defparam ram_block1a125.ram_block_type = "auto";

cycloneive_ram_block ram_block1a93(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[93]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a93_PORTBDATAOUT_bus));
defparam ram_block1a93.clk1_output_clock_enable = "ena1";
defparam ram_block1a93.data_interleave_offset_in_bits = 1;
defparam ram_block1a93.data_interleave_width_in_bits = 1;
defparam ram_block1a93.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a93.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a93.operation_mode = "dual_port";
defparam ram_block1a93.port_a_address_clear = "none";
defparam ram_block1a93.port_a_address_width = 3;
defparam ram_block1a93.port_a_data_out_clear = "none";
defparam ram_block1a93.port_a_data_out_clock = "none";
defparam ram_block1a93.port_a_data_width = 1;
defparam ram_block1a93.port_a_first_address = 0;
defparam ram_block1a93.port_a_first_bit_number = 93;
defparam ram_block1a93.port_a_last_address = 7;
defparam ram_block1a93.port_a_logical_ram_depth = 8;
defparam ram_block1a93.port_a_logical_ram_width = 258;
defparam ram_block1a93.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a93.port_b_address_clear = "none";
defparam ram_block1a93.port_b_address_clock = "clock1";
defparam ram_block1a93.port_b_address_width = 3;
defparam ram_block1a93.port_b_data_out_clear = "none";
defparam ram_block1a93.port_b_data_out_clock = "clock1";
defparam ram_block1a93.port_b_data_width = 1;
defparam ram_block1a93.port_b_first_address = 0;
defparam ram_block1a93.port_b_first_bit_number = 93;
defparam ram_block1a93.port_b_last_address = 7;
defparam ram_block1a93.port_b_logical_ram_depth = 8;
defparam ram_block1a93.port_b_logical_ram_width = 258;
defparam ram_block1a93.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a93.port_b_read_enable_clock = "clock1";
defparam ram_block1a93.ram_block_type = "auto";

cycloneive_ram_block ram_block1a77(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[77]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a77_PORTBDATAOUT_bus));
defparam ram_block1a77.clk1_output_clock_enable = "ena1";
defparam ram_block1a77.data_interleave_offset_in_bits = 1;
defparam ram_block1a77.data_interleave_width_in_bits = 1;
defparam ram_block1a77.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a77.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a77.operation_mode = "dual_port";
defparam ram_block1a77.port_a_address_clear = "none";
defparam ram_block1a77.port_a_address_width = 3;
defparam ram_block1a77.port_a_data_out_clear = "none";
defparam ram_block1a77.port_a_data_out_clock = "none";
defparam ram_block1a77.port_a_data_width = 1;
defparam ram_block1a77.port_a_first_address = 0;
defparam ram_block1a77.port_a_first_bit_number = 77;
defparam ram_block1a77.port_a_last_address = 7;
defparam ram_block1a77.port_a_logical_ram_depth = 8;
defparam ram_block1a77.port_a_logical_ram_width = 258;
defparam ram_block1a77.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a77.port_b_address_clear = "none";
defparam ram_block1a77.port_b_address_clock = "clock1";
defparam ram_block1a77.port_b_address_width = 3;
defparam ram_block1a77.port_b_data_out_clear = "none";
defparam ram_block1a77.port_b_data_out_clock = "clock1";
defparam ram_block1a77.port_b_data_width = 1;
defparam ram_block1a77.port_b_first_address = 0;
defparam ram_block1a77.port_b_first_bit_number = 77;
defparam ram_block1a77.port_b_last_address = 7;
defparam ram_block1a77.port_b_logical_ram_depth = 8;
defparam ram_block1a77.port_b_logical_ram_width = 258;
defparam ram_block1a77.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a77.port_b_read_enable_clock = "clock1";
defparam ram_block1a77.ram_block_type = "auto";

cycloneive_ram_block ram_block1a237(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[237]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a237_PORTBDATAOUT_bus));
defparam ram_block1a237.clk1_output_clock_enable = "ena1";
defparam ram_block1a237.data_interleave_offset_in_bits = 1;
defparam ram_block1a237.data_interleave_width_in_bits = 1;
defparam ram_block1a237.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a237.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a237.operation_mode = "dual_port";
defparam ram_block1a237.port_a_address_clear = "none";
defparam ram_block1a237.port_a_address_width = 3;
defparam ram_block1a237.port_a_data_out_clear = "none";
defparam ram_block1a237.port_a_data_out_clock = "none";
defparam ram_block1a237.port_a_data_width = 1;
defparam ram_block1a237.port_a_first_address = 0;
defparam ram_block1a237.port_a_first_bit_number = 237;
defparam ram_block1a237.port_a_last_address = 7;
defparam ram_block1a237.port_a_logical_ram_depth = 8;
defparam ram_block1a237.port_a_logical_ram_width = 258;
defparam ram_block1a237.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a237.port_b_address_clear = "none";
defparam ram_block1a237.port_b_address_clock = "clock1";
defparam ram_block1a237.port_b_address_width = 3;
defparam ram_block1a237.port_b_data_out_clear = "none";
defparam ram_block1a237.port_b_data_out_clock = "clock1";
defparam ram_block1a237.port_b_data_width = 1;
defparam ram_block1a237.port_b_first_address = 0;
defparam ram_block1a237.port_b_first_bit_number = 237;
defparam ram_block1a237.port_b_last_address = 7;
defparam ram_block1a237.port_b_logical_ram_depth = 8;
defparam ram_block1a237.port_b_logical_ram_width = 258;
defparam ram_block1a237.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a237.port_b_read_enable_clock = "clock1";
defparam ram_block1a237.ram_block_type = "auto";

cycloneive_ram_block ram_block1a253(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[253]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a253_PORTBDATAOUT_bus));
defparam ram_block1a253.clk1_output_clock_enable = "ena1";
defparam ram_block1a253.data_interleave_offset_in_bits = 1;
defparam ram_block1a253.data_interleave_width_in_bits = 1;
defparam ram_block1a253.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a253.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a253.operation_mode = "dual_port";
defparam ram_block1a253.port_a_address_clear = "none";
defparam ram_block1a253.port_a_address_width = 3;
defparam ram_block1a253.port_a_data_out_clear = "none";
defparam ram_block1a253.port_a_data_out_clock = "none";
defparam ram_block1a253.port_a_data_width = 1;
defparam ram_block1a253.port_a_first_address = 0;
defparam ram_block1a253.port_a_first_bit_number = 253;
defparam ram_block1a253.port_a_last_address = 7;
defparam ram_block1a253.port_a_logical_ram_depth = 8;
defparam ram_block1a253.port_a_logical_ram_width = 258;
defparam ram_block1a253.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a253.port_b_address_clear = "none";
defparam ram_block1a253.port_b_address_clock = "clock1";
defparam ram_block1a253.port_b_address_width = 3;
defparam ram_block1a253.port_b_data_out_clear = "none";
defparam ram_block1a253.port_b_data_out_clock = "clock1";
defparam ram_block1a253.port_b_data_width = 1;
defparam ram_block1a253.port_b_first_address = 0;
defparam ram_block1a253.port_b_first_bit_number = 253;
defparam ram_block1a253.port_b_last_address = 7;
defparam ram_block1a253.port_b_logical_ram_depth = 8;
defparam ram_block1a253.port_b_logical_ram_width = 258;
defparam ram_block1a253.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a253.port_b_read_enable_clock = "clock1";
defparam ram_block1a253.ram_block_type = "auto";

cycloneive_ram_block ram_block1a221(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[221]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a221_PORTBDATAOUT_bus));
defparam ram_block1a221.clk1_output_clock_enable = "ena1";
defparam ram_block1a221.data_interleave_offset_in_bits = 1;
defparam ram_block1a221.data_interleave_width_in_bits = 1;
defparam ram_block1a221.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a221.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a221.operation_mode = "dual_port";
defparam ram_block1a221.port_a_address_clear = "none";
defparam ram_block1a221.port_a_address_width = 3;
defparam ram_block1a221.port_a_data_out_clear = "none";
defparam ram_block1a221.port_a_data_out_clock = "none";
defparam ram_block1a221.port_a_data_width = 1;
defparam ram_block1a221.port_a_first_address = 0;
defparam ram_block1a221.port_a_first_bit_number = 221;
defparam ram_block1a221.port_a_last_address = 7;
defparam ram_block1a221.port_a_logical_ram_depth = 8;
defparam ram_block1a221.port_a_logical_ram_width = 258;
defparam ram_block1a221.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a221.port_b_address_clear = "none";
defparam ram_block1a221.port_b_address_clock = "clock1";
defparam ram_block1a221.port_b_address_width = 3;
defparam ram_block1a221.port_b_data_out_clear = "none";
defparam ram_block1a221.port_b_data_out_clock = "clock1";
defparam ram_block1a221.port_b_data_width = 1;
defparam ram_block1a221.port_b_first_address = 0;
defparam ram_block1a221.port_b_first_bit_number = 221;
defparam ram_block1a221.port_b_last_address = 7;
defparam ram_block1a221.port_b_logical_ram_depth = 8;
defparam ram_block1a221.port_b_logical_ram_width = 258;
defparam ram_block1a221.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a221.port_b_read_enable_clock = "clock1";
defparam ram_block1a221.ram_block_type = "auto";

cycloneive_ram_block ram_block1a205(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[205]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a205_PORTBDATAOUT_bus));
defparam ram_block1a205.clk1_output_clock_enable = "ena1";
defparam ram_block1a205.data_interleave_offset_in_bits = 1;
defparam ram_block1a205.data_interleave_width_in_bits = 1;
defparam ram_block1a205.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a205.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a205.operation_mode = "dual_port";
defparam ram_block1a205.port_a_address_clear = "none";
defparam ram_block1a205.port_a_address_width = 3;
defparam ram_block1a205.port_a_data_out_clear = "none";
defparam ram_block1a205.port_a_data_out_clock = "none";
defparam ram_block1a205.port_a_data_width = 1;
defparam ram_block1a205.port_a_first_address = 0;
defparam ram_block1a205.port_a_first_bit_number = 205;
defparam ram_block1a205.port_a_last_address = 7;
defparam ram_block1a205.port_a_logical_ram_depth = 8;
defparam ram_block1a205.port_a_logical_ram_width = 258;
defparam ram_block1a205.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a205.port_b_address_clear = "none";
defparam ram_block1a205.port_b_address_clock = "clock1";
defparam ram_block1a205.port_b_address_width = 3;
defparam ram_block1a205.port_b_data_out_clear = "none";
defparam ram_block1a205.port_b_data_out_clock = "clock1";
defparam ram_block1a205.port_b_data_width = 1;
defparam ram_block1a205.port_b_first_address = 0;
defparam ram_block1a205.port_b_first_bit_number = 205;
defparam ram_block1a205.port_b_last_address = 7;
defparam ram_block1a205.port_b_logical_ram_depth = 8;
defparam ram_block1a205.port_b_logical_ram_width = 258;
defparam ram_block1a205.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a205.port_b_read_enable_clock = "clock1";
defparam ram_block1a205.ram_block_type = "auto";

cycloneive_ram_block ram_block1a45(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[45]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a45_PORTBDATAOUT_bus));
defparam ram_block1a45.clk1_output_clock_enable = "ena1";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a45.operation_mode = "dual_port";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 3;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "none";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 0;
defparam ram_block1a45.port_a_first_bit_number = 45;
defparam ram_block1a45.port_a_last_address = 7;
defparam ram_block1a45.port_a_logical_ram_depth = 8;
defparam ram_block1a45.port_a_logical_ram_width = 258;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a45.port_b_address_clear = "none";
defparam ram_block1a45.port_b_address_clock = "clock1";
defparam ram_block1a45.port_b_address_width = 3;
defparam ram_block1a45.port_b_data_out_clear = "none";
defparam ram_block1a45.port_b_data_out_clock = "clock1";
defparam ram_block1a45.port_b_data_width = 1;
defparam ram_block1a45.port_b_first_address = 0;
defparam ram_block1a45.port_b_first_bit_number = 45;
defparam ram_block1a45.port_b_last_address = 7;
defparam ram_block1a45.port_b_logical_ram_depth = 8;
defparam ram_block1a45.port_b_logical_ram_width = 258;
defparam ram_block1a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a45.port_b_read_enable_clock = "clock1";
defparam ram_block1a45.ram_block_type = "auto";

cycloneive_ram_block ram_block1a61(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[61]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a61_PORTBDATAOUT_bus));
defparam ram_block1a61.clk1_output_clock_enable = "ena1";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a61.operation_mode = "dual_port";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 3;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "none";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 0;
defparam ram_block1a61.port_a_first_bit_number = 61;
defparam ram_block1a61.port_a_last_address = 7;
defparam ram_block1a61.port_a_logical_ram_depth = 8;
defparam ram_block1a61.port_a_logical_ram_width = 258;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a61.port_b_address_clear = "none";
defparam ram_block1a61.port_b_address_clock = "clock1";
defparam ram_block1a61.port_b_address_width = 3;
defparam ram_block1a61.port_b_data_out_clear = "none";
defparam ram_block1a61.port_b_data_out_clock = "clock1";
defparam ram_block1a61.port_b_data_width = 1;
defparam ram_block1a61.port_b_first_address = 0;
defparam ram_block1a61.port_b_first_bit_number = 61;
defparam ram_block1a61.port_b_last_address = 7;
defparam ram_block1a61.port_b_logical_ram_depth = 8;
defparam ram_block1a61.port_b_logical_ram_width = 258;
defparam ram_block1a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a61.port_b_read_enable_clock = "clock1";
defparam ram_block1a61.ram_block_type = "auto";

cycloneive_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk1_output_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 3;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 7;
defparam ram_block1a29.port_a_logical_ram_depth = 8;
defparam ram_block1a29.port_a_logical_ram_width = 258;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 3;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "clock1";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 7;
defparam ram_block1a29.port_b_logical_ram_depth = 8;
defparam ram_block1a29.port_b_logical_ram_width = 258;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 258;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 258;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a174(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[174]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a174_PORTBDATAOUT_bus));
defparam ram_block1a174.clk1_output_clock_enable = "ena1";
defparam ram_block1a174.data_interleave_offset_in_bits = 1;
defparam ram_block1a174.data_interleave_width_in_bits = 1;
defparam ram_block1a174.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a174.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a174.operation_mode = "dual_port";
defparam ram_block1a174.port_a_address_clear = "none";
defparam ram_block1a174.port_a_address_width = 3;
defparam ram_block1a174.port_a_data_out_clear = "none";
defparam ram_block1a174.port_a_data_out_clock = "none";
defparam ram_block1a174.port_a_data_width = 1;
defparam ram_block1a174.port_a_first_address = 0;
defparam ram_block1a174.port_a_first_bit_number = 174;
defparam ram_block1a174.port_a_last_address = 7;
defparam ram_block1a174.port_a_logical_ram_depth = 8;
defparam ram_block1a174.port_a_logical_ram_width = 258;
defparam ram_block1a174.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a174.port_b_address_clear = "none";
defparam ram_block1a174.port_b_address_clock = "clock1";
defparam ram_block1a174.port_b_address_width = 3;
defparam ram_block1a174.port_b_data_out_clear = "none";
defparam ram_block1a174.port_b_data_out_clock = "clock1";
defparam ram_block1a174.port_b_data_width = 1;
defparam ram_block1a174.port_b_first_address = 0;
defparam ram_block1a174.port_b_first_bit_number = 174;
defparam ram_block1a174.port_b_last_address = 7;
defparam ram_block1a174.port_b_logical_ram_depth = 8;
defparam ram_block1a174.port_b_logical_ram_width = 258;
defparam ram_block1a174.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a174.port_b_read_enable_clock = "clock1";
defparam ram_block1a174.ram_block_type = "auto";

cycloneive_ram_block ram_block1a110(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[110]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a110_PORTBDATAOUT_bus));
defparam ram_block1a110.clk1_output_clock_enable = "ena1";
defparam ram_block1a110.data_interleave_offset_in_bits = 1;
defparam ram_block1a110.data_interleave_width_in_bits = 1;
defparam ram_block1a110.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a110.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a110.operation_mode = "dual_port";
defparam ram_block1a110.port_a_address_clear = "none";
defparam ram_block1a110.port_a_address_width = 3;
defparam ram_block1a110.port_a_data_out_clear = "none";
defparam ram_block1a110.port_a_data_out_clock = "none";
defparam ram_block1a110.port_a_data_width = 1;
defparam ram_block1a110.port_a_first_address = 0;
defparam ram_block1a110.port_a_first_bit_number = 110;
defparam ram_block1a110.port_a_last_address = 7;
defparam ram_block1a110.port_a_logical_ram_depth = 8;
defparam ram_block1a110.port_a_logical_ram_width = 258;
defparam ram_block1a110.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a110.port_b_address_clear = "none";
defparam ram_block1a110.port_b_address_clock = "clock1";
defparam ram_block1a110.port_b_address_width = 3;
defparam ram_block1a110.port_b_data_out_clear = "none";
defparam ram_block1a110.port_b_data_out_clock = "clock1";
defparam ram_block1a110.port_b_data_width = 1;
defparam ram_block1a110.port_b_first_address = 0;
defparam ram_block1a110.port_b_first_bit_number = 110;
defparam ram_block1a110.port_b_last_address = 7;
defparam ram_block1a110.port_b_logical_ram_depth = 8;
defparam ram_block1a110.port_b_logical_ram_width = 258;
defparam ram_block1a110.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a110.port_b_read_enable_clock = "clock1";
defparam ram_block1a110.ram_block_type = "auto";

cycloneive_ram_block ram_block1a238(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[238]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a238_PORTBDATAOUT_bus));
defparam ram_block1a238.clk1_output_clock_enable = "ena1";
defparam ram_block1a238.data_interleave_offset_in_bits = 1;
defparam ram_block1a238.data_interleave_width_in_bits = 1;
defparam ram_block1a238.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a238.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a238.operation_mode = "dual_port";
defparam ram_block1a238.port_a_address_clear = "none";
defparam ram_block1a238.port_a_address_width = 3;
defparam ram_block1a238.port_a_data_out_clear = "none";
defparam ram_block1a238.port_a_data_out_clock = "none";
defparam ram_block1a238.port_a_data_width = 1;
defparam ram_block1a238.port_a_first_address = 0;
defparam ram_block1a238.port_a_first_bit_number = 238;
defparam ram_block1a238.port_a_last_address = 7;
defparam ram_block1a238.port_a_logical_ram_depth = 8;
defparam ram_block1a238.port_a_logical_ram_width = 258;
defparam ram_block1a238.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a238.port_b_address_clear = "none";
defparam ram_block1a238.port_b_address_clock = "clock1";
defparam ram_block1a238.port_b_address_width = 3;
defparam ram_block1a238.port_b_data_out_clear = "none";
defparam ram_block1a238.port_b_data_out_clock = "clock1";
defparam ram_block1a238.port_b_data_width = 1;
defparam ram_block1a238.port_b_first_address = 0;
defparam ram_block1a238.port_b_first_bit_number = 238;
defparam ram_block1a238.port_b_last_address = 7;
defparam ram_block1a238.port_b_logical_ram_depth = 8;
defparam ram_block1a238.port_b_logical_ram_width = 258;
defparam ram_block1a238.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a238.port_b_read_enable_clock = "clock1";
defparam ram_block1a238.ram_block_type = "auto";

cycloneive_ram_block ram_block1a46(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[46]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a46_PORTBDATAOUT_bus));
defparam ram_block1a46.clk1_output_clock_enable = "ena1";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a46.operation_mode = "dual_port";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 3;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "none";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 0;
defparam ram_block1a46.port_a_first_bit_number = 46;
defparam ram_block1a46.port_a_last_address = 7;
defparam ram_block1a46.port_a_logical_ram_depth = 8;
defparam ram_block1a46.port_a_logical_ram_width = 258;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a46.port_b_address_clear = "none";
defparam ram_block1a46.port_b_address_clock = "clock1";
defparam ram_block1a46.port_b_address_width = 3;
defparam ram_block1a46.port_b_data_out_clear = "none";
defparam ram_block1a46.port_b_data_out_clock = "clock1";
defparam ram_block1a46.port_b_data_width = 1;
defparam ram_block1a46.port_b_first_address = 0;
defparam ram_block1a46.port_b_first_bit_number = 46;
defparam ram_block1a46.port_b_last_address = 7;
defparam ram_block1a46.port_b_logical_ram_depth = 8;
defparam ram_block1a46.port_b_logical_ram_width = 258;
defparam ram_block1a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a46.port_b_read_enable_clock = "clock1";
defparam ram_block1a46.ram_block_type = "auto";

cycloneive_ram_block ram_block1a190(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[190]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a190_PORTBDATAOUT_bus));
defparam ram_block1a190.clk1_output_clock_enable = "ena1";
defparam ram_block1a190.data_interleave_offset_in_bits = 1;
defparam ram_block1a190.data_interleave_width_in_bits = 1;
defparam ram_block1a190.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a190.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a190.operation_mode = "dual_port";
defparam ram_block1a190.port_a_address_clear = "none";
defparam ram_block1a190.port_a_address_width = 3;
defparam ram_block1a190.port_a_data_out_clear = "none";
defparam ram_block1a190.port_a_data_out_clock = "none";
defparam ram_block1a190.port_a_data_width = 1;
defparam ram_block1a190.port_a_first_address = 0;
defparam ram_block1a190.port_a_first_bit_number = 190;
defparam ram_block1a190.port_a_last_address = 7;
defparam ram_block1a190.port_a_logical_ram_depth = 8;
defparam ram_block1a190.port_a_logical_ram_width = 258;
defparam ram_block1a190.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a190.port_b_address_clear = "none";
defparam ram_block1a190.port_b_address_clock = "clock1";
defparam ram_block1a190.port_b_address_width = 3;
defparam ram_block1a190.port_b_data_out_clear = "none";
defparam ram_block1a190.port_b_data_out_clock = "clock1";
defparam ram_block1a190.port_b_data_width = 1;
defparam ram_block1a190.port_b_first_address = 0;
defparam ram_block1a190.port_b_first_bit_number = 190;
defparam ram_block1a190.port_b_last_address = 7;
defparam ram_block1a190.port_b_logical_ram_depth = 8;
defparam ram_block1a190.port_b_logical_ram_width = 258;
defparam ram_block1a190.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a190.port_b_read_enable_clock = "clock1";
defparam ram_block1a190.ram_block_type = "auto";

cycloneive_ram_block ram_block1a126(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[126]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a126_PORTBDATAOUT_bus));
defparam ram_block1a126.clk1_output_clock_enable = "ena1";
defparam ram_block1a126.data_interleave_offset_in_bits = 1;
defparam ram_block1a126.data_interleave_width_in_bits = 1;
defparam ram_block1a126.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a126.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a126.operation_mode = "dual_port";
defparam ram_block1a126.port_a_address_clear = "none";
defparam ram_block1a126.port_a_address_width = 3;
defparam ram_block1a126.port_a_data_out_clear = "none";
defparam ram_block1a126.port_a_data_out_clock = "none";
defparam ram_block1a126.port_a_data_width = 1;
defparam ram_block1a126.port_a_first_address = 0;
defparam ram_block1a126.port_a_first_bit_number = 126;
defparam ram_block1a126.port_a_last_address = 7;
defparam ram_block1a126.port_a_logical_ram_depth = 8;
defparam ram_block1a126.port_a_logical_ram_width = 258;
defparam ram_block1a126.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a126.port_b_address_clear = "none";
defparam ram_block1a126.port_b_address_clock = "clock1";
defparam ram_block1a126.port_b_address_width = 3;
defparam ram_block1a126.port_b_data_out_clear = "none";
defparam ram_block1a126.port_b_data_out_clock = "clock1";
defparam ram_block1a126.port_b_data_width = 1;
defparam ram_block1a126.port_b_first_address = 0;
defparam ram_block1a126.port_b_first_bit_number = 126;
defparam ram_block1a126.port_b_last_address = 7;
defparam ram_block1a126.port_b_logical_ram_depth = 8;
defparam ram_block1a126.port_b_logical_ram_width = 258;
defparam ram_block1a126.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a126.port_b_read_enable_clock = "clock1";
defparam ram_block1a126.ram_block_type = "auto";

cycloneive_ram_block ram_block1a254(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[254]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a254_PORTBDATAOUT_bus));
defparam ram_block1a254.clk1_output_clock_enable = "ena1";
defparam ram_block1a254.data_interleave_offset_in_bits = 1;
defparam ram_block1a254.data_interleave_width_in_bits = 1;
defparam ram_block1a254.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a254.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a254.operation_mode = "dual_port";
defparam ram_block1a254.port_a_address_clear = "none";
defparam ram_block1a254.port_a_address_width = 3;
defparam ram_block1a254.port_a_data_out_clear = "none";
defparam ram_block1a254.port_a_data_out_clock = "none";
defparam ram_block1a254.port_a_data_width = 1;
defparam ram_block1a254.port_a_first_address = 0;
defparam ram_block1a254.port_a_first_bit_number = 254;
defparam ram_block1a254.port_a_last_address = 7;
defparam ram_block1a254.port_a_logical_ram_depth = 8;
defparam ram_block1a254.port_a_logical_ram_width = 258;
defparam ram_block1a254.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a254.port_b_address_clear = "none";
defparam ram_block1a254.port_b_address_clock = "clock1";
defparam ram_block1a254.port_b_address_width = 3;
defparam ram_block1a254.port_b_data_out_clear = "none";
defparam ram_block1a254.port_b_data_out_clock = "clock1";
defparam ram_block1a254.port_b_data_width = 1;
defparam ram_block1a254.port_b_first_address = 0;
defparam ram_block1a254.port_b_first_bit_number = 254;
defparam ram_block1a254.port_b_last_address = 7;
defparam ram_block1a254.port_b_logical_ram_depth = 8;
defparam ram_block1a254.port_b_logical_ram_width = 258;
defparam ram_block1a254.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a254.port_b_read_enable_clock = "clock1";
defparam ram_block1a254.ram_block_type = "auto";

cycloneive_ram_block ram_block1a62(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[62]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a62_PORTBDATAOUT_bus));
defparam ram_block1a62.clk1_output_clock_enable = "ena1";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a62.operation_mode = "dual_port";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 3;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "none";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 0;
defparam ram_block1a62.port_a_first_bit_number = 62;
defparam ram_block1a62.port_a_last_address = 7;
defparam ram_block1a62.port_a_logical_ram_depth = 8;
defparam ram_block1a62.port_a_logical_ram_width = 258;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a62.port_b_address_clear = "none";
defparam ram_block1a62.port_b_address_clock = "clock1";
defparam ram_block1a62.port_b_address_width = 3;
defparam ram_block1a62.port_b_data_out_clear = "none";
defparam ram_block1a62.port_b_data_out_clock = "clock1";
defparam ram_block1a62.port_b_data_width = 1;
defparam ram_block1a62.port_b_first_address = 0;
defparam ram_block1a62.port_b_first_bit_number = 62;
defparam ram_block1a62.port_b_last_address = 7;
defparam ram_block1a62.port_b_logical_ram_depth = 8;
defparam ram_block1a62.port_b_logical_ram_width = 258;
defparam ram_block1a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a62.port_b_read_enable_clock = "clock1";
defparam ram_block1a62.ram_block_type = "auto";

cycloneive_ram_block ram_block1a94(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[94]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a94_PORTBDATAOUT_bus));
defparam ram_block1a94.clk1_output_clock_enable = "ena1";
defparam ram_block1a94.data_interleave_offset_in_bits = 1;
defparam ram_block1a94.data_interleave_width_in_bits = 1;
defparam ram_block1a94.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a94.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a94.operation_mode = "dual_port";
defparam ram_block1a94.port_a_address_clear = "none";
defparam ram_block1a94.port_a_address_width = 3;
defparam ram_block1a94.port_a_data_out_clear = "none";
defparam ram_block1a94.port_a_data_out_clock = "none";
defparam ram_block1a94.port_a_data_width = 1;
defparam ram_block1a94.port_a_first_address = 0;
defparam ram_block1a94.port_a_first_bit_number = 94;
defparam ram_block1a94.port_a_last_address = 7;
defparam ram_block1a94.port_a_logical_ram_depth = 8;
defparam ram_block1a94.port_a_logical_ram_width = 258;
defparam ram_block1a94.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a94.port_b_address_clear = "none";
defparam ram_block1a94.port_b_address_clock = "clock1";
defparam ram_block1a94.port_b_address_width = 3;
defparam ram_block1a94.port_b_data_out_clear = "none";
defparam ram_block1a94.port_b_data_out_clock = "clock1";
defparam ram_block1a94.port_b_data_width = 1;
defparam ram_block1a94.port_b_first_address = 0;
defparam ram_block1a94.port_b_first_bit_number = 94;
defparam ram_block1a94.port_b_last_address = 7;
defparam ram_block1a94.port_b_logical_ram_depth = 8;
defparam ram_block1a94.port_b_logical_ram_width = 258;
defparam ram_block1a94.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a94.port_b_read_enable_clock = "clock1";
defparam ram_block1a94.ram_block_type = "auto";

cycloneive_ram_block ram_block1a158(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[158]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a158_PORTBDATAOUT_bus));
defparam ram_block1a158.clk1_output_clock_enable = "ena1";
defparam ram_block1a158.data_interleave_offset_in_bits = 1;
defparam ram_block1a158.data_interleave_width_in_bits = 1;
defparam ram_block1a158.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a158.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a158.operation_mode = "dual_port";
defparam ram_block1a158.port_a_address_clear = "none";
defparam ram_block1a158.port_a_address_width = 3;
defparam ram_block1a158.port_a_data_out_clear = "none";
defparam ram_block1a158.port_a_data_out_clock = "none";
defparam ram_block1a158.port_a_data_width = 1;
defparam ram_block1a158.port_a_first_address = 0;
defparam ram_block1a158.port_a_first_bit_number = 158;
defparam ram_block1a158.port_a_last_address = 7;
defparam ram_block1a158.port_a_logical_ram_depth = 8;
defparam ram_block1a158.port_a_logical_ram_width = 258;
defparam ram_block1a158.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a158.port_b_address_clear = "none";
defparam ram_block1a158.port_b_address_clock = "clock1";
defparam ram_block1a158.port_b_address_width = 3;
defparam ram_block1a158.port_b_data_out_clear = "none";
defparam ram_block1a158.port_b_data_out_clock = "clock1";
defparam ram_block1a158.port_b_data_width = 1;
defparam ram_block1a158.port_b_first_address = 0;
defparam ram_block1a158.port_b_first_bit_number = 158;
defparam ram_block1a158.port_b_last_address = 7;
defparam ram_block1a158.port_b_logical_ram_depth = 8;
defparam ram_block1a158.port_b_logical_ram_width = 258;
defparam ram_block1a158.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a158.port_b_read_enable_clock = "clock1";
defparam ram_block1a158.ram_block_type = "auto";

cycloneive_ram_block ram_block1a222(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[222]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a222_PORTBDATAOUT_bus));
defparam ram_block1a222.clk1_output_clock_enable = "ena1";
defparam ram_block1a222.data_interleave_offset_in_bits = 1;
defparam ram_block1a222.data_interleave_width_in_bits = 1;
defparam ram_block1a222.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a222.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a222.operation_mode = "dual_port";
defparam ram_block1a222.port_a_address_clear = "none";
defparam ram_block1a222.port_a_address_width = 3;
defparam ram_block1a222.port_a_data_out_clear = "none";
defparam ram_block1a222.port_a_data_out_clock = "none";
defparam ram_block1a222.port_a_data_width = 1;
defparam ram_block1a222.port_a_first_address = 0;
defparam ram_block1a222.port_a_first_bit_number = 222;
defparam ram_block1a222.port_a_last_address = 7;
defparam ram_block1a222.port_a_logical_ram_depth = 8;
defparam ram_block1a222.port_a_logical_ram_width = 258;
defparam ram_block1a222.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a222.port_b_address_clear = "none";
defparam ram_block1a222.port_b_address_clock = "clock1";
defparam ram_block1a222.port_b_address_width = 3;
defparam ram_block1a222.port_b_data_out_clear = "none";
defparam ram_block1a222.port_b_data_out_clock = "clock1";
defparam ram_block1a222.port_b_data_width = 1;
defparam ram_block1a222.port_b_first_address = 0;
defparam ram_block1a222.port_b_first_bit_number = 222;
defparam ram_block1a222.port_b_last_address = 7;
defparam ram_block1a222.port_b_logical_ram_depth = 8;
defparam ram_block1a222.port_b_logical_ram_width = 258;
defparam ram_block1a222.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a222.port_b_read_enable_clock = "clock1";
defparam ram_block1a222.ram_block_type = "auto";

cycloneive_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk1_output_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 3;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 7;
defparam ram_block1a30.port_a_logical_ram_depth = 8;
defparam ram_block1a30.port_a_logical_ram_width = 258;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 3;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "clock1";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 7;
defparam ram_block1a30.port_b_logical_ram_depth = 8;
defparam ram_block1a30.port_b_logical_ram_width = 258;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cycloneive_ram_block ram_block1a78(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[78]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a78_PORTBDATAOUT_bus));
defparam ram_block1a78.clk1_output_clock_enable = "ena1";
defparam ram_block1a78.data_interleave_offset_in_bits = 1;
defparam ram_block1a78.data_interleave_width_in_bits = 1;
defparam ram_block1a78.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a78.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a78.operation_mode = "dual_port";
defparam ram_block1a78.port_a_address_clear = "none";
defparam ram_block1a78.port_a_address_width = 3;
defparam ram_block1a78.port_a_data_out_clear = "none";
defparam ram_block1a78.port_a_data_out_clock = "none";
defparam ram_block1a78.port_a_data_width = 1;
defparam ram_block1a78.port_a_first_address = 0;
defparam ram_block1a78.port_a_first_bit_number = 78;
defparam ram_block1a78.port_a_last_address = 7;
defparam ram_block1a78.port_a_logical_ram_depth = 8;
defparam ram_block1a78.port_a_logical_ram_width = 258;
defparam ram_block1a78.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a78.port_b_address_clear = "none";
defparam ram_block1a78.port_b_address_clock = "clock1";
defparam ram_block1a78.port_b_address_width = 3;
defparam ram_block1a78.port_b_data_out_clear = "none";
defparam ram_block1a78.port_b_data_out_clock = "clock1";
defparam ram_block1a78.port_b_data_width = 1;
defparam ram_block1a78.port_b_first_address = 0;
defparam ram_block1a78.port_b_first_bit_number = 78;
defparam ram_block1a78.port_b_last_address = 7;
defparam ram_block1a78.port_b_logical_ram_depth = 8;
defparam ram_block1a78.port_b_logical_ram_width = 258;
defparam ram_block1a78.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a78.port_b_read_enable_clock = "clock1";
defparam ram_block1a78.ram_block_type = "auto";

cycloneive_ram_block ram_block1a142(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[142]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a142_PORTBDATAOUT_bus));
defparam ram_block1a142.clk1_output_clock_enable = "ena1";
defparam ram_block1a142.data_interleave_offset_in_bits = 1;
defparam ram_block1a142.data_interleave_width_in_bits = 1;
defparam ram_block1a142.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a142.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a142.operation_mode = "dual_port";
defparam ram_block1a142.port_a_address_clear = "none";
defparam ram_block1a142.port_a_address_width = 3;
defparam ram_block1a142.port_a_data_out_clear = "none";
defparam ram_block1a142.port_a_data_out_clock = "none";
defparam ram_block1a142.port_a_data_width = 1;
defparam ram_block1a142.port_a_first_address = 0;
defparam ram_block1a142.port_a_first_bit_number = 142;
defparam ram_block1a142.port_a_last_address = 7;
defparam ram_block1a142.port_a_logical_ram_depth = 8;
defparam ram_block1a142.port_a_logical_ram_width = 258;
defparam ram_block1a142.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a142.port_b_address_clear = "none";
defparam ram_block1a142.port_b_address_clock = "clock1";
defparam ram_block1a142.port_b_address_width = 3;
defparam ram_block1a142.port_b_data_out_clear = "none";
defparam ram_block1a142.port_b_data_out_clock = "clock1";
defparam ram_block1a142.port_b_data_width = 1;
defparam ram_block1a142.port_b_first_address = 0;
defparam ram_block1a142.port_b_first_bit_number = 142;
defparam ram_block1a142.port_b_last_address = 7;
defparam ram_block1a142.port_b_logical_ram_depth = 8;
defparam ram_block1a142.port_b_logical_ram_width = 258;
defparam ram_block1a142.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a142.port_b_read_enable_clock = "clock1";
defparam ram_block1a142.ram_block_type = "auto";

cycloneive_ram_block ram_block1a206(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[206]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a206_PORTBDATAOUT_bus));
defparam ram_block1a206.clk1_output_clock_enable = "ena1";
defparam ram_block1a206.data_interleave_offset_in_bits = 1;
defparam ram_block1a206.data_interleave_width_in_bits = 1;
defparam ram_block1a206.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a206.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a206.operation_mode = "dual_port";
defparam ram_block1a206.port_a_address_clear = "none";
defparam ram_block1a206.port_a_address_width = 3;
defparam ram_block1a206.port_a_data_out_clear = "none";
defparam ram_block1a206.port_a_data_out_clock = "none";
defparam ram_block1a206.port_a_data_width = 1;
defparam ram_block1a206.port_a_first_address = 0;
defparam ram_block1a206.port_a_first_bit_number = 206;
defparam ram_block1a206.port_a_last_address = 7;
defparam ram_block1a206.port_a_logical_ram_depth = 8;
defparam ram_block1a206.port_a_logical_ram_width = 258;
defparam ram_block1a206.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a206.port_b_address_clear = "none";
defparam ram_block1a206.port_b_address_clock = "clock1";
defparam ram_block1a206.port_b_address_width = 3;
defparam ram_block1a206.port_b_data_out_clear = "none";
defparam ram_block1a206.port_b_data_out_clock = "clock1";
defparam ram_block1a206.port_b_data_width = 1;
defparam ram_block1a206.port_b_first_address = 0;
defparam ram_block1a206.port_b_first_bit_number = 206;
defparam ram_block1a206.port_b_last_address = 7;
defparam ram_block1a206.port_b_logical_ram_depth = 8;
defparam ram_block1a206.port_b_logical_ram_width = 258;
defparam ram_block1a206.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a206.port_b_read_enable_clock = "clock1";
defparam ram_block1a206.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 258;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 258;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a111(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[111]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a111_PORTBDATAOUT_bus));
defparam ram_block1a111.clk1_output_clock_enable = "ena1";
defparam ram_block1a111.data_interleave_offset_in_bits = 1;
defparam ram_block1a111.data_interleave_width_in_bits = 1;
defparam ram_block1a111.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a111.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a111.operation_mode = "dual_port";
defparam ram_block1a111.port_a_address_clear = "none";
defparam ram_block1a111.port_a_address_width = 3;
defparam ram_block1a111.port_a_data_out_clear = "none";
defparam ram_block1a111.port_a_data_out_clock = "none";
defparam ram_block1a111.port_a_data_width = 1;
defparam ram_block1a111.port_a_first_address = 0;
defparam ram_block1a111.port_a_first_bit_number = 111;
defparam ram_block1a111.port_a_last_address = 7;
defparam ram_block1a111.port_a_logical_ram_depth = 8;
defparam ram_block1a111.port_a_logical_ram_width = 258;
defparam ram_block1a111.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a111.port_b_address_clear = "none";
defparam ram_block1a111.port_b_address_clock = "clock1";
defparam ram_block1a111.port_b_address_width = 3;
defparam ram_block1a111.port_b_data_out_clear = "none";
defparam ram_block1a111.port_b_data_out_clock = "clock1";
defparam ram_block1a111.port_b_data_width = 1;
defparam ram_block1a111.port_b_first_address = 0;
defparam ram_block1a111.port_b_first_bit_number = 111;
defparam ram_block1a111.port_b_last_address = 7;
defparam ram_block1a111.port_b_logical_ram_depth = 8;
defparam ram_block1a111.port_b_logical_ram_width = 258;
defparam ram_block1a111.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a111.port_b_read_enable_clock = "clock1";
defparam ram_block1a111.ram_block_type = "auto";

cycloneive_ram_block ram_block1a127(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[127]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a127_PORTBDATAOUT_bus));
defparam ram_block1a127.clk1_output_clock_enable = "ena1";
defparam ram_block1a127.data_interleave_offset_in_bits = 1;
defparam ram_block1a127.data_interleave_width_in_bits = 1;
defparam ram_block1a127.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a127.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a127.operation_mode = "dual_port";
defparam ram_block1a127.port_a_address_clear = "none";
defparam ram_block1a127.port_a_address_width = 3;
defparam ram_block1a127.port_a_data_out_clear = "none";
defparam ram_block1a127.port_a_data_out_clock = "none";
defparam ram_block1a127.port_a_data_width = 1;
defparam ram_block1a127.port_a_first_address = 0;
defparam ram_block1a127.port_a_first_bit_number = 127;
defparam ram_block1a127.port_a_last_address = 7;
defparam ram_block1a127.port_a_logical_ram_depth = 8;
defparam ram_block1a127.port_a_logical_ram_width = 258;
defparam ram_block1a127.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a127.port_b_address_clear = "none";
defparam ram_block1a127.port_b_address_clock = "clock1";
defparam ram_block1a127.port_b_address_width = 3;
defparam ram_block1a127.port_b_data_out_clear = "none";
defparam ram_block1a127.port_b_data_out_clock = "clock1";
defparam ram_block1a127.port_b_data_width = 1;
defparam ram_block1a127.port_b_first_address = 0;
defparam ram_block1a127.port_b_first_bit_number = 127;
defparam ram_block1a127.port_b_last_address = 7;
defparam ram_block1a127.port_b_logical_ram_depth = 8;
defparam ram_block1a127.port_b_logical_ram_width = 258;
defparam ram_block1a127.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a127.port_b_read_enable_clock = "clock1";
defparam ram_block1a127.ram_block_type = "auto";

cycloneive_ram_block ram_block1a95(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[95]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a95_PORTBDATAOUT_bus));
defparam ram_block1a95.clk1_output_clock_enable = "ena1";
defparam ram_block1a95.data_interleave_offset_in_bits = 1;
defparam ram_block1a95.data_interleave_width_in_bits = 1;
defparam ram_block1a95.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a95.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a95.operation_mode = "dual_port";
defparam ram_block1a95.port_a_address_clear = "none";
defparam ram_block1a95.port_a_address_width = 3;
defparam ram_block1a95.port_a_data_out_clear = "none";
defparam ram_block1a95.port_a_data_out_clock = "none";
defparam ram_block1a95.port_a_data_width = 1;
defparam ram_block1a95.port_a_first_address = 0;
defparam ram_block1a95.port_a_first_bit_number = 95;
defparam ram_block1a95.port_a_last_address = 7;
defparam ram_block1a95.port_a_logical_ram_depth = 8;
defparam ram_block1a95.port_a_logical_ram_width = 258;
defparam ram_block1a95.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a95.port_b_address_clear = "none";
defparam ram_block1a95.port_b_address_clock = "clock1";
defparam ram_block1a95.port_b_address_width = 3;
defparam ram_block1a95.port_b_data_out_clear = "none";
defparam ram_block1a95.port_b_data_out_clock = "clock1";
defparam ram_block1a95.port_b_data_width = 1;
defparam ram_block1a95.port_b_first_address = 0;
defparam ram_block1a95.port_b_first_bit_number = 95;
defparam ram_block1a95.port_b_last_address = 7;
defparam ram_block1a95.port_b_logical_ram_depth = 8;
defparam ram_block1a95.port_b_logical_ram_width = 258;
defparam ram_block1a95.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a95.port_b_read_enable_clock = "clock1";
defparam ram_block1a95.ram_block_type = "auto";

cycloneive_ram_block ram_block1a79(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[79]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a79_PORTBDATAOUT_bus));
defparam ram_block1a79.clk1_output_clock_enable = "ena1";
defparam ram_block1a79.data_interleave_offset_in_bits = 1;
defparam ram_block1a79.data_interleave_width_in_bits = 1;
defparam ram_block1a79.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a79.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a79.operation_mode = "dual_port";
defparam ram_block1a79.port_a_address_clear = "none";
defparam ram_block1a79.port_a_address_width = 3;
defparam ram_block1a79.port_a_data_out_clear = "none";
defparam ram_block1a79.port_a_data_out_clock = "none";
defparam ram_block1a79.port_a_data_width = 1;
defparam ram_block1a79.port_a_first_address = 0;
defparam ram_block1a79.port_a_first_bit_number = 79;
defparam ram_block1a79.port_a_last_address = 7;
defparam ram_block1a79.port_a_logical_ram_depth = 8;
defparam ram_block1a79.port_a_logical_ram_width = 258;
defparam ram_block1a79.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a79.port_b_address_clear = "none";
defparam ram_block1a79.port_b_address_clock = "clock1";
defparam ram_block1a79.port_b_address_width = 3;
defparam ram_block1a79.port_b_data_out_clear = "none";
defparam ram_block1a79.port_b_data_out_clock = "clock1";
defparam ram_block1a79.port_b_data_width = 1;
defparam ram_block1a79.port_b_first_address = 0;
defparam ram_block1a79.port_b_first_bit_number = 79;
defparam ram_block1a79.port_b_last_address = 7;
defparam ram_block1a79.port_b_logical_ram_depth = 8;
defparam ram_block1a79.port_b_logical_ram_width = 258;
defparam ram_block1a79.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a79.port_b_read_enable_clock = "clock1";
defparam ram_block1a79.ram_block_type = "auto";

cycloneive_ram_block ram_block1a175(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[175]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a175_PORTBDATAOUT_bus));
defparam ram_block1a175.clk1_output_clock_enable = "ena1";
defparam ram_block1a175.data_interleave_offset_in_bits = 1;
defparam ram_block1a175.data_interleave_width_in_bits = 1;
defparam ram_block1a175.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a175.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a175.operation_mode = "dual_port";
defparam ram_block1a175.port_a_address_clear = "none";
defparam ram_block1a175.port_a_address_width = 3;
defparam ram_block1a175.port_a_data_out_clear = "none";
defparam ram_block1a175.port_a_data_out_clock = "none";
defparam ram_block1a175.port_a_data_width = 1;
defparam ram_block1a175.port_a_first_address = 0;
defparam ram_block1a175.port_a_first_bit_number = 175;
defparam ram_block1a175.port_a_last_address = 7;
defparam ram_block1a175.port_a_logical_ram_depth = 8;
defparam ram_block1a175.port_a_logical_ram_width = 258;
defparam ram_block1a175.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a175.port_b_address_clear = "none";
defparam ram_block1a175.port_b_address_clock = "clock1";
defparam ram_block1a175.port_b_address_width = 3;
defparam ram_block1a175.port_b_data_out_clear = "none";
defparam ram_block1a175.port_b_data_out_clock = "clock1";
defparam ram_block1a175.port_b_data_width = 1;
defparam ram_block1a175.port_b_first_address = 0;
defparam ram_block1a175.port_b_first_bit_number = 175;
defparam ram_block1a175.port_b_last_address = 7;
defparam ram_block1a175.port_b_logical_ram_depth = 8;
defparam ram_block1a175.port_b_logical_ram_width = 258;
defparam ram_block1a175.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a175.port_b_read_enable_clock = "clock1";
defparam ram_block1a175.ram_block_type = "auto";

cycloneive_ram_block ram_block1a191(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[191]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a191_PORTBDATAOUT_bus));
defparam ram_block1a191.clk1_output_clock_enable = "ena1";
defparam ram_block1a191.data_interleave_offset_in_bits = 1;
defparam ram_block1a191.data_interleave_width_in_bits = 1;
defparam ram_block1a191.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a191.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a191.operation_mode = "dual_port";
defparam ram_block1a191.port_a_address_clear = "none";
defparam ram_block1a191.port_a_address_width = 3;
defparam ram_block1a191.port_a_data_out_clear = "none";
defparam ram_block1a191.port_a_data_out_clock = "none";
defparam ram_block1a191.port_a_data_width = 1;
defparam ram_block1a191.port_a_first_address = 0;
defparam ram_block1a191.port_a_first_bit_number = 191;
defparam ram_block1a191.port_a_last_address = 7;
defparam ram_block1a191.port_a_logical_ram_depth = 8;
defparam ram_block1a191.port_a_logical_ram_width = 258;
defparam ram_block1a191.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a191.port_b_address_clear = "none";
defparam ram_block1a191.port_b_address_clock = "clock1";
defparam ram_block1a191.port_b_address_width = 3;
defparam ram_block1a191.port_b_data_out_clear = "none";
defparam ram_block1a191.port_b_data_out_clock = "clock1";
defparam ram_block1a191.port_b_data_width = 1;
defparam ram_block1a191.port_b_first_address = 0;
defparam ram_block1a191.port_b_first_bit_number = 191;
defparam ram_block1a191.port_b_last_address = 7;
defparam ram_block1a191.port_b_logical_ram_depth = 8;
defparam ram_block1a191.port_b_logical_ram_width = 258;
defparam ram_block1a191.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a191.port_b_read_enable_clock = "clock1";
defparam ram_block1a191.ram_block_type = "auto";

cycloneive_ram_block ram_block1a159(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[159]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a159_PORTBDATAOUT_bus));
defparam ram_block1a159.clk1_output_clock_enable = "ena1";
defparam ram_block1a159.data_interleave_offset_in_bits = 1;
defparam ram_block1a159.data_interleave_width_in_bits = 1;
defparam ram_block1a159.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a159.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a159.operation_mode = "dual_port";
defparam ram_block1a159.port_a_address_clear = "none";
defparam ram_block1a159.port_a_address_width = 3;
defparam ram_block1a159.port_a_data_out_clear = "none";
defparam ram_block1a159.port_a_data_out_clock = "none";
defparam ram_block1a159.port_a_data_width = 1;
defparam ram_block1a159.port_a_first_address = 0;
defparam ram_block1a159.port_a_first_bit_number = 159;
defparam ram_block1a159.port_a_last_address = 7;
defparam ram_block1a159.port_a_logical_ram_depth = 8;
defparam ram_block1a159.port_a_logical_ram_width = 258;
defparam ram_block1a159.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a159.port_b_address_clear = "none";
defparam ram_block1a159.port_b_address_clock = "clock1";
defparam ram_block1a159.port_b_address_width = 3;
defparam ram_block1a159.port_b_data_out_clear = "none";
defparam ram_block1a159.port_b_data_out_clock = "clock1";
defparam ram_block1a159.port_b_data_width = 1;
defparam ram_block1a159.port_b_first_address = 0;
defparam ram_block1a159.port_b_first_bit_number = 159;
defparam ram_block1a159.port_b_last_address = 7;
defparam ram_block1a159.port_b_logical_ram_depth = 8;
defparam ram_block1a159.port_b_logical_ram_width = 258;
defparam ram_block1a159.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a159.port_b_read_enable_clock = "clock1";
defparam ram_block1a159.ram_block_type = "auto";

cycloneive_ram_block ram_block1a143(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[143]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a143_PORTBDATAOUT_bus));
defparam ram_block1a143.clk1_output_clock_enable = "ena1";
defparam ram_block1a143.data_interleave_offset_in_bits = 1;
defparam ram_block1a143.data_interleave_width_in_bits = 1;
defparam ram_block1a143.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a143.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a143.operation_mode = "dual_port";
defparam ram_block1a143.port_a_address_clear = "none";
defparam ram_block1a143.port_a_address_width = 3;
defparam ram_block1a143.port_a_data_out_clear = "none";
defparam ram_block1a143.port_a_data_out_clock = "none";
defparam ram_block1a143.port_a_data_width = 1;
defparam ram_block1a143.port_a_first_address = 0;
defparam ram_block1a143.port_a_first_bit_number = 143;
defparam ram_block1a143.port_a_last_address = 7;
defparam ram_block1a143.port_a_logical_ram_depth = 8;
defparam ram_block1a143.port_a_logical_ram_width = 258;
defparam ram_block1a143.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a143.port_b_address_clear = "none";
defparam ram_block1a143.port_b_address_clock = "clock1";
defparam ram_block1a143.port_b_address_width = 3;
defparam ram_block1a143.port_b_data_out_clear = "none";
defparam ram_block1a143.port_b_data_out_clock = "clock1";
defparam ram_block1a143.port_b_data_width = 1;
defparam ram_block1a143.port_b_first_address = 0;
defparam ram_block1a143.port_b_first_bit_number = 143;
defparam ram_block1a143.port_b_last_address = 7;
defparam ram_block1a143.port_b_logical_ram_depth = 8;
defparam ram_block1a143.port_b_logical_ram_width = 258;
defparam ram_block1a143.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a143.port_b_read_enable_clock = "clock1";
defparam ram_block1a143.ram_block_type = "auto";

cycloneive_ram_block ram_block1a239(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[239]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a239_PORTBDATAOUT_bus));
defparam ram_block1a239.clk1_output_clock_enable = "ena1";
defparam ram_block1a239.data_interleave_offset_in_bits = 1;
defparam ram_block1a239.data_interleave_width_in_bits = 1;
defparam ram_block1a239.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a239.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a239.operation_mode = "dual_port";
defparam ram_block1a239.port_a_address_clear = "none";
defparam ram_block1a239.port_a_address_width = 3;
defparam ram_block1a239.port_a_data_out_clear = "none";
defparam ram_block1a239.port_a_data_out_clock = "none";
defparam ram_block1a239.port_a_data_width = 1;
defparam ram_block1a239.port_a_first_address = 0;
defparam ram_block1a239.port_a_first_bit_number = 239;
defparam ram_block1a239.port_a_last_address = 7;
defparam ram_block1a239.port_a_logical_ram_depth = 8;
defparam ram_block1a239.port_a_logical_ram_width = 258;
defparam ram_block1a239.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a239.port_b_address_clear = "none";
defparam ram_block1a239.port_b_address_clock = "clock1";
defparam ram_block1a239.port_b_address_width = 3;
defparam ram_block1a239.port_b_data_out_clear = "none";
defparam ram_block1a239.port_b_data_out_clock = "clock1";
defparam ram_block1a239.port_b_data_width = 1;
defparam ram_block1a239.port_b_first_address = 0;
defparam ram_block1a239.port_b_first_bit_number = 239;
defparam ram_block1a239.port_b_last_address = 7;
defparam ram_block1a239.port_b_logical_ram_depth = 8;
defparam ram_block1a239.port_b_logical_ram_width = 258;
defparam ram_block1a239.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a239.port_b_read_enable_clock = "clock1";
defparam ram_block1a239.ram_block_type = "auto";

cycloneive_ram_block ram_block1a255(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[255]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a255_PORTBDATAOUT_bus));
defparam ram_block1a255.clk1_output_clock_enable = "ena1";
defparam ram_block1a255.data_interleave_offset_in_bits = 1;
defparam ram_block1a255.data_interleave_width_in_bits = 1;
defparam ram_block1a255.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a255.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a255.operation_mode = "dual_port";
defparam ram_block1a255.port_a_address_clear = "none";
defparam ram_block1a255.port_a_address_width = 3;
defparam ram_block1a255.port_a_data_out_clear = "none";
defparam ram_block1a255.port_a_data_out_clock = "none";
defparam ram_block1a255.port_a_data_width = 1;
defparam ram_block1a255.port_a_first_address = 0;
defparam ram_block1a255.port_a_first_bit_number = 255;
defparam ram_block1a255.port_a_last_address = 7;
defparam ram_block1a255.port_a_logical_ram_depth = 8;
defparam ram_block1a255.port_a_logical_ram_width = 258;
defparam ram_block1a255.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a255.port_b_address_clear = "none";
defparam ram_block1a255.port_b_address_clock = "clock1";
defparam ram_block1a255.port_b_address_width = 3;
defparam ram_block1a255.port_b_data_out_clear = "none";
defparam ram_block1a255.port_b_data_out_clock = "clock1";
defparam ram_block1a255.port_b_data_width = 1;
defparam ram_block1a255.port_b_first_address = 0;
defparam ram_block1a255.port_b_first_bit_number = 255;
defparam ram_block1a255.port_b_last_address = 7;
defparam ram_block1a255.port_b_logical_ram_depth = 8;
defparam ram_block1a255.port_b_logical_ram_width = 258;
defparam ram_block1a255.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a255.port_b_read_enable_clock = "clock1";
defparam ram_block1a255.ram_block_type = "auto";

cycloneive_ram_block ram_block1a223(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[223]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a223_PORTBDATAOUT_bus));
defparam ram_block1a223.clk1_output_clock_enable = "ena1";
defparam ram_block1a223.data_interleave_offset_in_bits = 1;
defparam ram_block1a223.data_interleave_width_in_bits = 1;
defparam ram_block1a223.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a223.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a223.operation_mode = "dual_port";
defparam ram_block1a223.port_a_address_clear = "none";
defparam ram_block1a223.port_a_address_width = 3;
defparam ram_block1a223.port_a_data_out_clear = "none";
defparam ram_block1a223.port_a_data_out_clock = "none";
defparam ram_block1a223.port_a_data_width = 1;
defparam ram_block1a223.port_a_first_address = 0;
defparam ram_block1a223.port_a_first_bit_number = 223;
defparam ram_block1a223.port_a_last_address = 7;
defparam ram_block1a223.port_a_logical_ram_depth = 8;
defparam ram_block1a223.port_a_logical_ram_width = 258;
defparam ram_block1a223.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a223.port_b_address_clear = "none";
defparam ram_block1a223.port_b_address_clock = "clock1";
defparam ram_block1a223.port_b_address_width = 3;
defparam ram_block1a223.port_b_data_out_clear = "none";
defparam ram_block1a223.port_b_data_out_clock = "clock1";
defparam ram_block1a223.port_b_data_width = 1;
defparam ram_block1a223.port_b_first_address = 0;
defparam ram_block1a223.port_b_first_bit_number = 223;
defparam ram_block1a223.port_b_last_address = 7;
defparam ram_block1a223.port_b_logical_ram_depth = 8;
defparam ram_block1a223.port_b_logical_ram_width = 258;
defparam ram_block1a223.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a223.port_b_read_enable_clock = "clock1";
defparam ram_block1a223.ram_block_type = "auto";

cycloneive_ram_block ram_block1a207(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[207]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a207_PORTBDATAOUT_bus));
defparam ram_block1a207.clk1_output_clock_enable = "ena1";
defparam ram_block1a207.data_interleave_offset_in_bits = 1;
defparam ram_block1a207.data_interleave_width_in_bits = 1;
defparam ram_block1a207.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a207.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a207.operation_mode = "dual_port";
defparam ram_block1a207.port_a_address_clear = "none";
defparam ram_block1a207.port_a_address_width = 3;
defparam ram_block1a207.port_a_data_out_clear = "none";
defparam ram_block1a207.port_a_data_out_clock = "none";
defparam ram_block1a207.port_a_data_width = 1;
defparam ram_block1a207.port_a_first_address = 0;
defparam ram_block1a207.port_a_first_bit_number = 207;
defparam ram_block1a207.port_a_last_address = 7;
defparam ram_block1a207.port_a_logical_ram_depth = 8;
defparam ram_block1a207.port_a_logical_ram_width = 258;
defparam ram_block1a207.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a207.port_b_address_clear = "none";
defparam ram_block1a207.port_b_address_clock = "clock1";
defparam ram_block1a207.port_b_address_width = 3;
defparam ram_block1a207.port_b_data_out_clear = "none";
defparam ram_block1a207.port_b_data_out_clock = "clock1";
defparam ram_block1a207.port_b_data_width = 1;
defparam ram_block1a207.port_b_first_address = 0;
defparam ram_block1a207.port_b_first_bit_number = 207;
defparam ram_block1a207.port_b_last_address = 7;
defparam ram_block1a207.port_b_logical_ram_depth = 8;
defparam ram_block1a207.port_b_logical_ram_width = 258;
defparam ram_block1a207.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a207.port_b_read_enable_clock = "clock1";
defparam ram_block1a207.ram_block_type = "auto";

cycloneive_ram_block ram_block1a47(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[47]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a47_PORTBDATAOUT_bus));
defparam ram_block1a47.clk1_output_clock_enable = "ena1";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a47.operation_mode = "dual_port";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 3;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "none";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 0;
defparam ram_block1a47.port_a_first_bit_number = 47;
defparam ram_block1a47.port_a_last_address = 7;
defparam ram_block1a47.port_a_logical_ram_depth = 8;
defparam ram_block1a47.port_a_logical_ram_width = 258;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a47.port_b_address_clear = "none";
defparam ram_block1a47.port_b_address_clock = "clock1";
defparam ram_block1a47.port_b_address_width = 3;
defparam ram_block1a47.port_b_data_out_clear = "none";
defparam ram_block1a47.port_b_data_out_clock = "clock1";
defparam ram_block1a47.port_b_data_width = 1;
defparam ram_block1a47.port_b_first_address = 0;
defparam ram_block1a47.port_b_first_bit_number = 47;
defparam ram_block1a47.port_b_last_address = 7;
defparam ram_block1a47.port_b_logical_ram_depth = 8;
defparam ram_block1a47.port_b_logical_ram_width = 258;
defparam ram_block1a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a47.port_b_read_enable_clock = "clock1";
defparam ram_block1a47.ram_block_type = "auto";

cycloneive_ram_block ram_block1a63(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[63]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a63_PORTBDATAOUT_bus));
defparam ram_block1a63.clk1_output_clock_enable = "ena1";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a63.operation_mode = "dual_port";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 3;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "none";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 0;
defparam ram_block1a63.port_a_first_bit_number = 63;
defparam ram_block1a63.port_a_last_address = 7;
defparam ram_block1a63.port_a_logical_ram_depth = 8;
defparam ram_block1a63.port_a_logical_ram_width = 258;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a63.port_b_address_clear = "none";
defparam ram_block1a63.port_b_address_clock = "clock1";
defparam ram_block1a63.port_b_address_width = 3;
defparam ram_block1a63.port_b_data_out_clear = "none";
defparam ram_block1a63.port_b_data_out_clock = "clock1";
defparam ram_block1a63.port_b_data_width = 1;
defparam ram_block1a63.port_b_first_address = 0;
defparam ram_block1a63.port_b_first_bit_number = 63;
defparam ram_block1a63.port_b_last_address = 7;
defparam ram_block1a63.port_b_logical_ram_depth = 8;
defparam ram_block1a63.port_b_logical_ram_width = 258;
defparam ram_block1a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a63.port_b_read_enable_clock = "clock1";
defparam ram_block1a63.ram_block_type = "auto";

cycloneive_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk1_output_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 3;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 7;
defparam ram_block1a31.port_a_logical_ram_depth = 8;
defparam ram_block1a31.port_a_logical_ram_width = 258;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 3;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "clock1";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 7;
defparam ram_block1a31.port_b_logical_ram_depth = 8;
defparam ram_block1a31.port_b_logical_ram_width = 258;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_6h71:auto_generated|a_dpfifo_nmv:dpfifo|altsyncram_1bh1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 258;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 258;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

endmodule

module CIC_cntr_8a7 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	valid_rreq,
	updown,
	GND_port,
	clock,
	in_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	valid_rreq;
input 	updown;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~2_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~2 (
	.dataa(in_valid),
	.datab(full_dff),
	.datac(valid_rreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'h96FF;
defparam \_~2 .sum_lutc_input = "datac";

endmodule

module CIC_cntr_r9b (
	counter_reg_bit_0,
	counter_reg_bit_1,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout());
defparam counter_comb_bita1.lut_mask = 16'h5A5A;
defparam counter_comb_bita1.sum_lutc_input = "cin";

endmodule

module CIC_cntr_s9b (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	GND_port,
	clock,
	in_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(in_valid),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module CIC_auk_dspip_avalon_streaming_source (
	at_source_data,
	source_valid_s1,
	at_source_channel,
	dffe_af,
	state_0,
	data,
	stall_reg,
	dout_valid,
	data_count,
	GND_port,
	clk,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[15:0] at_source_data;
output 	source_valid_s1;
output 	[3:0] at_source_channel;
output 	dffe_af;
input 	state_0;
input 	[15:0] data;
input 	stall_reg;
input 	dout_valid;
input 	[3:0] data_count;
input 	GND_port;
input 	clk;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \source_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \source_valid_s_process~0_combout ;


CIC_scfifo_18 source_FIFO(
	.q({q_unconnected_wire_257,q_unconnected_wire_256,q_unconnected_wire_255,q_unconnected_wire_254,q_unconnected_wire_253,q_unconnected_wire_252,q_unconnected_wire_251,q_unconnected_wire_250,q_unconnected_wire_249,q_unconnected_wire_248,q_unconnected_wire_247,
q_unconnected_wire_246,q_unconnected_wire_245,q_unconnected_wire_244,q_unconnected_wire_243,q_unconnected_wire_242,q_unconnected_wire_241,q_unconnected_wire_240,q_unconnected_wire_239,q_unconnected_wire_238,q_unconnected_wire_237,q_unconnected_wire_236,
q_unconnected_wire_235,q_unconnected_wire_234,q_unconnected_wire_233,q_unconnected_wire_232,q_unconnected_wire_231,q_unconnected_wire_230,q_unconnected_wire_229,q_unconnected_wire_228,q_unconnected_wire_227,q_unconnected_wire_226,q_unconnected_wire_225,
q_unconnected_wire_224,q_unconnected_wire_223,q_unconnected_wire_222,q_unconnected_wire_221,q_unconnected_wire_220,q_unconnected_wire_219,q_unconnected_wire_218,q_unconnected_wire_217,q_unconnected_wire_216,q_unconnected_wire_215,q_unconnected_wire_214,
q_unconnected_wire_213,q_unconnected_wire_212,q_unconnected_wire_211,q_unconnected_wire_210,q_unconnected_wire_209,q_unconnected_wire_208,q_unconnected_wire_207,q_unconnected_wire_206,q_unconnected_wire_205,q_unconnected_wire_204,q_unconnected_wire_203,
q_unconnected_wire_202,q_unconnected_wire_201,q_unconnected_wire_200,q_unconnected_wire_199,q_unconnected_wire_198,q_unconnected_wire_197,q_unconnected_wire_196,q_unconnected_wire_195,q_unconnected_wire_194,q_unconnected_wire_193,q_unconnected_wire_192,
q_unconnected_wire_191,q_unconnected_wire_190,q_unconnected_wire_189,q_unconnected_wire_188,q_unconnected_wire_187,q_unconnected_wire_186,q_unconnected_wire_185,q_unconnected_wire_184,q_unconnected_wire_183,q_unconnected_wire_182,q_unconnected_wire_181,
q_unconnected_wire_180,q_unconnected_wire_179,q_unconnected_wire_178,q_unconnected_wire_177,q_unconnected_wire_176,q_unconnected_wire_175,q_unconnected_wire_174,q_unconnected_wire_173,q_unconnected_wire_172,q_unconnected_wire_171,q_unconnected_wire_170,
q_unconnected_wire_169,q_unconnected_wire_168,q_unconnected_wire_167,q_unconnected_wire_166,q_unconnected_wire_165,q_unconnected_wire_164,q_unconnected_wire_163,q_unconnected_wire_162,q_unconnected_wire_161,q_unconnected_wire_160,q_unconnected_wire_159,
q_unconnected_wire_158,q_unconnected_wire_157,q_unconnected_wire_156,q_unconnected_wire_155,q_unconnected_wire_154,q_unconnected_wire_153,q_unconnected_wire_152,q_unconnected_wire_151,q_unconnected_wire_150,q_unconnected_wire_149,q_unconnected_wire_148,
q_unconnected_wire_147,q_unconnected_wire_146,q_unconnected_wire_145,q_unconnected_wire_144,q_unconnected_wire_143,q_unconnected_wire_142,q_unconnected_wire_141,q_unconnected_wire_140,q_unconnected_wire_139,q_unconnected_wire_138,q_unconnected_wire_137,
q_unconnected_wire_136,q_unconnected_wire_135,q_unconnected_wire_134,q_unconnected_wire_133,q_unconnected_wire_132,q_unconnected_wire_131,q_unconnected_wire_130,q_unconnected_wire_129,q_unconnected_wire_128,q_unconnected_wire_127,q_unconnected_wire_126,
q_unconnected_wire_125,q_unconnected_wire_124,q_unconnected_wire_123,q_unconnected_wire_122,q_unconnected_wire_121,q_unconnected_wire_120,q_unconnected_wire_119,q_unconnected_wire_118,q_unconnected_wire_117,q_unconnected_wire_116,q_unconnected_wire_115,
q_unconnected_wire_114,q_unconnected_wire_113,q_unconnected_wire_112,q_unconnected_wire_111,q_unconnected_wire_110,q_unconnected_wire_109,q_unconnected_wire_108,q_unconnected_wire_107,q_unconnected_wire_106,q_unconnected_wire_105,q_unconnected_wire_104,
q_unconnected_wire_103,q_unconnected_wire_102,q_unconnected_wire_101,q_unconnected_wire_100,q_unconnected_wire_99,q_unconnected_wire_98,q_unconnected_wire_97,q_unconnected_wire_96,q_unconnected_wire_95,q_unconnected_wire_94,q_unconnected_wire_93,q_unconnected_wire_92,
q_unconnected_wire_91,q_unconnected_wire_90,q_unconnected_wire_89,q_unconnected_wire_88,q_unconnected_wire_87,q_unconnected_wire_86,q_unconnected_wire_85,q_unconnected_wire_84,q_unconnected_wire_83,q_unconnected_wire_82,q_unconnected_wire_81,q_unconnected_wire_80,
q_unconnected_wire_79,q_unconnected_wire_78,q_unconnected_wire_77,q_unconnected_wire_76,q_unconnected_wire_75,q_unconnected_wire_74,q_unconnected_wire_73,q_unconnected_wire_72,q_unconnected_wire_71,q_unconnected_wire_70,q_unconnected_wire_69,q_unconnected_wire_68,
q_unconnected_wire_67,q_unconnected_wire_66,q_unconnected_wire_65,q_unconnected_wire_64,q_unconnected_wire_63,q_unconnected_wire_62,q_unconnected_wire_61,q_unconnected_wire_60,q_unconnected_wire_59,q_unconnected_wire_58,q_unconnected_wire_57,q_unconnected_wire_56,
q_unconnected_wire_55,q_unconnected_wire_54,q_unconnected_wire_53,q_unconnected_wire_52,q_unconnected_wire_51,q_unconnected_wire_50,q_unconnected_wire_49,q_unconnected_wire_48,q_unconnected_wire_47,q_unconnected_wire_46,q_unconnected_wire_45,q_unconnected_wire_44,
q_unconnected_wire_43,q_unconnected_wire_42,q_unconnected_wire_41,q_unconnected_wire_40,q_unconnected_wire_39,q_unconnected_wire_38,q_unconnected_wire_37,q_unconnected_wire_36,q_unconnected_wire_35,q_unconnected_wire_34,q_unconnected_wire_33,q_unconnected_wire_32,
q_unconnected_wire_31,q_unconnected_wire_30,q_unconnected_wire_29,q_unconnected_wire_28,q_unconnected_wire_27,q_unconnected_wire_26,q_unconnected_wire_25,q_unconnected_wire_24,q_unconnected_wire_23,q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,
at_source_channel[3],at_source_channel[2],at_source_channel[1],at_source_channel[0],at_source_data[15],at_source_data[14],at_source_data[13],at_source_data[12],at_source_data[11],at_source_data[10],at_source_data[9],at_source_data[8],at_source_data[7],at_source_data[6],at_source_data[5],at_source_data[4],at_source_data[3],
at_source_data[2],at_source_data[1],at_source_data[0]}),
	.source_valid_s(source_valid_s1),
	.dffe_af(dffe_af),
	.state_0(state_0),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_count[3],data_count[2],data_count[1],data_count[0],data[15],data[14],data[13],
data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid),
	.empty_dff(\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n),
	.out_ready(out_ready));

dffeas source_valid_s(
	.clk(clk),
	.d(\source_valid_s_process~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(source_valid_s1),
	.prn(vcc));
defparam source_valid_s.is_wysiwyg = "true";
defparam source_valid_s.power_up = "low";

cycloneive_lcell_comb \source_valid_s_process~0 (
	.dataa(out_ready),
	.datab(gnd),
	.datac(source_valid_s1),
	.datad(\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.cin(gnd),
	.combout(\source_valid_s_process~0_combout ),
	.cout());
defparam \source_valid_s_process~0 .lut_mask = 16'hFFF5;
defparam \source_valid_s_process~0 .sum_lutc_input = "datac";

endmodule

module CIC_scfifo_18 (
	q,
	source_valid_s,
	dffe_af,
	state_0,
	data,
	stall_reg,
	dout_valid,
	empty_dff,
	GND_port,
	clock,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[257:0] q;
input 	source_valid_s;
output 	dffe_af;
input 	state_0;
input 	[257:0] data;
input 	stall_reg;
input 	dout_valid;
output 	empty_dff;
input 	GND_port;
input 	clock;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



CIC_scfifo_6i71 auto_generated(
	.q({q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.source_valid_s(source_valid_s),
	.dffe_af1(dffe_af),
	.state_0(state_0),
	.data({data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid),
	.empty_dff(empty_dff),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n),
	.out_ready(out_ready));

endmodule

module CIC_scfifo_6i71 (
	q,
	source_valid_s,
	dffe_af1,
	state_0,
	data,
	stall_reg,
	dout_valid,
	empty_dff,
	GND_port,
	clock,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q;
input 	source_valid_s;
output 	dffe_af1;
input 	state_0;
input 	[19:0] data;
input 	stall_reg;
input 	dout_valid;
output 	empty_dff;
input 	GND_port;
input 	clock;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;
wire \dffe_af~2_combout ;
wire \dffe_af~3_combout ;


CIC_a_dpfifo_3qv dpfifo(
	.q({q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.source_valid_s(source_valid_s),
	.state_0(state_0),
	.data({data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_4(\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_0(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid),
	.empty_dff1(empty_dff),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n),
	.out_ready(out_ready));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

cycloneive_lcell_comb \dffe_af~0 (
	.dataa(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datac(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datad(\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.cin(gnd),
	.combout(\dffe_af~0_combout ),
	.cout());
defparam \dffe_af~0 .lut_mask = 16'hEFFF;
defparam \dffe_af~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe_af~1 (
	.dataa(stall_reg),
	.datab(dout_valid),
	.datac(state_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\dffe_af~1_combout ),
	.cout());
defparam \dffe_af~1 .lut_mask = 16'hFDFD;
defparam \dffe_af~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe_af~2 (
	.dataa(dffe_af1),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(source_valid_s),
	.datad(out_ready),
	.cin(gnd),
	.combout(\dffe_af~2_combout ),
	.cout());
defparam \dffe_af~2 .lut_mask = 16'h6996;
defparam \dffe_af~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dffe_af~3 (
	.dataa(\dffe_af~0_combout ),
	.datab(\dffe_af~1_combout ),
	.datac(dffe_af1),
	.datad(\dffe_af~2_combout ),
	.cin(gnd),
	.combout(\dffe_af~3_combout ),
	.cout());
defparam \dffe_af~3 .lut_mask = 16'hFDFE;
defparam \dffe_af~3 .sum_lutc_input = "datac";

endmodule

module CIC_a_dpfifo_3qv (
	q,
	source_valid_s,
	state_0,
	data,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_0,
	stall_reg,
	dout_valid,
	empty_dff1,
	GND_port,
	clock,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q;
input 	source_valid_s;
input 	state_0;
input 	[19:0] data;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
input 	stall_reg;
input 	dout_valid;
output 	empty_dff1;
input 	GND_port;
input 	clock;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;
wire \usedw_is_0_dff~q ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \full_dff~q ;
wire \valid_wreq~combout ;
wire \valid_rreq~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \empty_dff~1_combout ;


CIC_cntr_u9b_16 wr_ptr(
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(\valid_wreq~combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_aa7_16 usedw_counter(
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_0(counter_reg_bit_0),
	.updown(\valid_wreq~combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_cntr_t9b_16 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

CIC_altsyncram_5ah1 FIFOram(
	.q_b({q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock1(clock),
	.clock0(clock));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

cycloneive_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

cycloneive_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rd_ptr_lsb~1 (
	.dataa(empty_dff1),
	.datab(out_ready),
	.datac(source_valid_s),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

cycloneive_lcell_comb \_~2 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hBFFF;
defparam \_~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~3 (
	.dataa(\full_dff~q ),
	.datab(counter_reg_bit_4),
	.datac(\_~2_combout ),
	.datad(\valid_wreq~combout ),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFEFF;
defparam \_~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \_~4 (
	.dataa(empty_dff1),
	.datab(out_ready),
	.datac(source_valid_s),
	.datad(\_~3_combout ),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hFFF7;
defparam \_~4 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

cycloneive_lcell_comb valid_wreq(
	.dataa(\full_dff~q ),
	.datab(stall_reg),
	.datac(dout_valid),
	.datad(state_0),
	.cin(gnd),
	.combout(\valid_wreq~combout ),
	.cout());
defparam valid_wreq.lut_mask = 16'hEFFF;
defparam valid_wreq.sum_lutc_input = "datac";

cycloneive_lcell_comb \valid_rreq~0 (
	.dataa(empty_dff1),
	.datab(out_ready),
	.datac(gnd),
	.datad(source_valid_s),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~0 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'h7FFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~1 (
	.dataa(\valid_wreq~combout ),
	.datab(\valid_rreq~0_combout ),
	.datac(counter_reg_bit_1),
	.datad(\usedw_will_be_1~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\usedw_is_0_dff~q ),
	.datac(\valid_wreq~combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFB;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFEFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

cycloneive_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~combout ),
	.datac(\valid_rreq~0_combout ),
	.datad(\usedw_is_1_dff~q ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBEFF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hFEFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

endmodule

module CIC_altsyncram_5ah1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[19:0] q_b;
input 	[19:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

cycloneive_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 20;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 20;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cycloneive_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 20;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 20;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cycloneive_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 20;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 20;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cycloneive_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 20;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 20;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cycloneive_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 20;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 20;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cycloneive_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 20;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 20;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cycloneive_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 20;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 20;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cycloneive_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 20;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 20;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cycloneive_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 20;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 20;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cycloneive_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 20;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 20;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cycloneive_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 20;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 20;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cycloneive_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 20;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 20;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cycloneive_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 20;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 20;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cycloneive_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 20;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 20;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cycloneive_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 20;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 20;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cycloneive_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 20;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 20;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cycloneive_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 20;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 20;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cycloneive_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 20;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 20;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cycloneive_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 20;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 20;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cycloneive_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "CIC_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_6i71:auto_generated|a_dpfifo_3qv:dpfifo|altsyncram_5ah1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 20;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 20;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

endmodule

module CIC_cntr_aa7_16 (
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_0,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(updown),
	.datab(valid_rreq),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h66FF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module CIC_cntr_t9b_16 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module CIC_cntr_u9b_16 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

cycloneive_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

cycloneive_lcell_comb \_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(reset_n),
	.datad(valid_wreq),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h0FFF;
defparam \_~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

cycloneive_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule
