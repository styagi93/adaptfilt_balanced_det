��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[/�������]�4wE�tO�$�2s۰,v`['�@��J�S2w�2<��E�k��[{�>�FA�T� )���y�*�
3��Bm���&=�S6_��ɛ�gz�=v��P�������\[��]6	���8�����?'�U�
9����C���P�=K�	+55�xƦ����-m8j����
a�./Wc:�����Nd�6�T#�n�H �E�o����	V�7٦Mx^`�]�q5��f��&��"f�]��օ~��:��Ӯ-h㋅�ݢ��u��ؿ��L&��I�i�ȧ�c��q��m��8dD*;l�і?po�3W���I �J�湡�}6H	`� ���5�{�E@?+j3�6i*؇��P��=Z�Y%o�}� �M��<���;  s;1����������Q��uQ�.�.20l��(�MQͩf�b= ���r��s�zO#���I.�Q�&���������Uo��z2�e[=J�N�ěД�T�/�$�6Y3�6ʘ���p8��*�oPu�\_еh�~�+*r1�L�Ϊ	,��O#��� �~�f���,Yn��"n&9 �_��>n�03�$-���r�	eJ�nx��=�ϯ��&�TM�����úCڂ����&�?7ѹG�g�fn�L�����I���Nm@*# �F?��Ƥ�\�Q|��^�n1�Ve|�XQx�|�i�Zm�c����;)����V�
��<��)�q2���vǋĲ&��<OZ�ꍲT�P�R����J(�,g������J��8���YĂ�$�n�ϣU�O��b`(��=�I������S�G.� ���+�VFq[��Y�ƴin�n���x��� A֮i#��@��|#a��a��2b����V�DU��� g�l��7G�bdkq�M6.��C�Ӊ/�9Т�����R��U[�J�8�_�U��qߺ������\����W��
�C��</,
R^���	��3	J�J���6D��M���q�k�H�P@���������]t=Y0��ЏiT���k?@�=��t5�P/���^�vׯũ��q�(��aO�Ĳ�CA�N����Q�e0�VW�?I�T�!��H�\X�p�$?B
a�W.�0sb��)U���	�I	�l�Gx��<��0[z�%"*�)��wt���R�����q�_�	m}M�H�
�>g����#|h�y�t�2[�2���eQ�Ce��'�5^�E�w�˧�g|�a���u�ɝ+��E��2pB��wm���T�|�?I�=����>�UM�C�IA����>�Ԧ�U����Y,�ʓ��Q���cLN�I�, Ƴ����{}#Hd�W9��@<����������� ����x���y�A=�UZ�?��t=������_'����=��}���IԖ'�&3�38ͧT����Q,ɾ�4X��_���hBT)b��?��Ѭ�2F�ƺ�Nڇ5�?;��|����N�/���͋����|��Z��t�ѿ{7Ģe\[�F�ƩG{�i�j��� �Ж)u����%O[�>�&�hˇ�9�U�K`�F׌P�:�5�d��Wn���+wL`i��P���5]�v�^�Yޛb��� G��0B|�`���#d�I:�a=[�X�m��H/��`C|+���_öG\`%�c8D9x8��+^vKZ�$q4�. {5�n�J�.$hl���ȼ�V�3	�iYD  �s
�Vb�Kd�4Hu!���y�a�}��s齧�ʺ0ϱZH|Mr���83�i�ۮg���+�fm	o���i�=+��;u�#Y����1�aنy����(�E���N��!Y��K:2�E�6�,�m�P�6W���ߨ����F�"��ڡ(�����[/Q��}�f����*��ȃ���p$
nh[��]3mp�s'5�Z%�\q\(q�<��:t�'���q��2��.૳�J��
J��+�|�-2b�ۮ�07���ж��J�=ޙɓ	_G(��ʇ�1>$&���ZJ��
�a�`(��bWPN	���]�T����뇪��.����c��f^��V@S�s:h�p�O�R�+!N��qG�&�0��_�j� =�$��i;��yo�̍ٶn{�)���,²�f(��	\v��.�bM��g�W��*���!���?�:�x?S���,5�܏���O+�i��K;�	L	MG� C��,ӱA��:��q��D"~�Ǆkŗ��a��ϥ�E�b[w�'Pī����Z��~����28��C��n���ͽъ����Y�:������{Go�-����B?DQu$$��_�zoe�Wvi�~�8<��/�Ȉ.�6-�S�DڮT�����_�g����?0�ULD��Gj�S<����;/���
�3&HL�?v�ƛ뀐�}�7|�>R�����2P�����x��ϼa.��KA�	51�q��u0/��2�ۚZ��I����<R�����P�6��7�f����I3W"�m���~����x�F%�U-`�|�f\�{���H��F<G�j1|id�r���L`jvC�&Vm%
Pw�¬Z��x �"�E�u�=�m&�ǘB�W��J��i��1�w���
fZ
���:�0���:���L��T4Bv�_g�dT���Xl��z�^�`$h�O�!Q��X<�U5H7��߭B0ط�Hk��wA�w�nz쥶8��i�w'�`z�b�"g��Â5E҅�R�U�T�"E+��[ȋ�]���Du�`\t� )������Q�v��0#ƽ3�X����B6Ĝ�r���u�4,,I5#jYS�{�T'Y�X'�"�cG b:�`,|��*�ή�����<*d�V�'L�cˀ�A6-�]��-�l+�!i��a�%4c�P�Mk�hN?ja�n��L}DR�v��`d�U��.u6{��E'��,�3�a��b�R~j��q���w�ؕ��
B��/�]<�[p��%M�v��r�Ŷ���՞!c��*���c���r(�PQ�V��	m�H��K/@D�������%h�c��I�!�{���s��E�u�0#��2���~l&��)-��%����ώl�� ��sb�;�GT�p��A����jC���)�8NB?�=<\ (�O���Uh=l�װ��w�H�G�!��7�J4Q�bBM�C����`�;<�KG��s���UI��QRp�r� pX)l+�B""�f������x^V�]���v�7��$�KOj�_��@��}��i��s#�v�-�1^g���9s��]�;�\����h=��������M/й��Ѱ
�sY'��C|#�P
��
[}�u���ʂ������1 �'�X���쎓�W�T��!�տ+��[�DhaKo�a�kԉ�Wf��c�>��`4(�&�4�5Iq��4/%�BO�eD�{��3���U.$�G��]X�{�|\g�*��Y>��p3��;|��C��k[,H�͗w6���}91�M�i��LYϳ��TB��imL�p�@/�K�{�I.r5]�N�7�Ou�t��$2������!��bIW����&��'xO=�s�`|>B�B�����B�!���r�R��>R�N�/�d�0���yT;����p5��b�uꬊ�ܧ���a^�3�2ڀ�&��Ʌa������[ �4�k0���5/�^P�=����_�0"�34��/)�f���&�zO7g�5�u�Tn����H6`��P�;"�Ԛ�u�vN�P�"�n��%UF�D��(�PŃ��	F�t�,�� a7���I�vPX$��s�UD$M�/�^�c����b�h����R0�9�1��Wɸ�yޤ�췀i�"/�c�=)&<��W���7��|45��U�]"x��GC��� l��R_��<Mê_���L��c�^vtXtAYP���׮��\Z�烧��ǴUz�2�|u�bu�m�\��,n~\�R�R�p�O���i����q��B��S\��Iw�Z��8��p�}���];���|{~���of������\fm@`��8��a�g3������x���/m�̬�V�-�7�Nv��Q�	$x�r�br��ZX=�Y��t���̲�im�pr k��5�3y6�� p�2@��и>_�� �^�*B��,��F�E� �C ��#� ��:g]n%�����i� ٢?D���Th�����֪�ɖy�\ۯ@Ԝ���\���Zɬt%�r��%�CC���������EMU�lo�P`|o�u������q \2T�ё�.�`��ܯN�(\T,&�:D}s[�7�O�0�#춈S���a�=(��@%*���B+�Ҥ|fi����)��P��Q9�W���5v��K���P�|�;�$yxU�i	;`��=�u�V�0�窭)w����фz}Y直�x����ڒ]��������%%b��]��*N]`�����{���S	Awl��"#��a�
#e�OsyQ(:]��t��[����,��ƭ��K󷃡yDO�+�SV�:����'
�~z�ǎ�!A0j��%A -�7�K[�m�������.��<.��v"!e9�cf�����д&��DKD<?��P��w�W�Dɨ=`ZgV�b����A���X�:���s��t5p����,�~��K��E=�蠞�?ֆ�i���C���D]㘰;{q=��8�>㠩|#�JZ:�M�CN�G�_�Y�����Ye����O�����c�R��8/%+��pR��ѹ��t�*�>��x�L��eu{a�$�A���gL�o�����Q�R�g�ϭ��it�D��-<�`Z�|��U4uN�k'�F�{��E^ձK2K�tI℧>��h���hDF��{�)�<���
`�p�;m���{q\ Q�aI�W�!��y���_�����58����dh��>+����y��'<W�/K3�|���9X��5C��1�����f
�_��O�_� ��{Q0�0y��Ԣ�Z�Ԁd�*���O��C �����HV5�r���g��-�%�^�i�����R	�����9S1�,k�O'M�ވC"Ij����x�5��[�P��(-��K�k�ۼ�~�6�k��~F7�ݪ�K�W�� 4aw;��V�h�z��w��!nL�^���F�����ޥG��!#qu�����݆n}�����@��^�
�{� ΈF����� ;2��P�WKsis`��y`�����{]�� ,s�au�R�8�؏Ϊ}k8Fb��|6��hXW��9yIS�Mpc���9N� F��E�N1B���l5�C�,I{-���3��k.�*�
�@Tbx���kƨ��Yd��=K�0���.����l�7n�eL��ʡ�͆��NCMT��a4IM[V�%���
?��b1J�nS�s�|�+8w!��d��
�!�YA7�(c ���j��
#�Β}�ߙI��]
6B�)1�i�)?w���  ���\�}ዦn�#��7��D<����]e?f ��]| ��y��|��1����#�Gg�j3L#JP�-��E�3M!c�P`IC��:�o�ݑ,`��<b�dD�}�-����rs�SJ'�ְU#aG�^/��1��%��J  ��Q�,���&�զK�3�m�va6z���LoN*��{o��2��h����S��ӵ�_�z�2��db0�ǡ�a*�5�o�h���h1Y=�|}� qn��P~�Ͽ�U�69�V+G�3D�C�I�Y��x�!��ρ��'"^jR�RO2o�B𭔳%n鴽��c7���x~��gl�g��Ex�A��bWM�B��E��7�c���v3�at���R儬���2�9�ի�����Y#��J�԰��ϳ�)���O{4M���wk���H�������	 ���?E'(�ER.�J��+�W�!��g����P>i���
��òzI�8�B;|,�{�-�I�	>A��e�g`5c���Gm˻!CA������1qLv^�ɪ�|�C5jĉ�:��\�O���ܙ��F SO�;����U��-������8M�
i68"��D�-IR��9y�g�c���8�	?yV�)Z�p�N���@t1W�����N�,�*�
4��j�d��nz��ge���nE-�س�~t��ܝ��ävʋD�	�a[��)��$g9��T���oۢm��-��� eĎ�$��5��/�s��^��ffc�~i��2$6_�܁������5��$���j�wK�����0	�C��$��T���j��[��)�D�� w6�;	%����hn���>����Ġ��Pmk$��9���j�o<&*X�Xe��^�'"W�Aݟۭ�q	T�1} �JfK�#t	 �u�go`_���A31_�p�e�@Xs�q��㚽y�Kk�֡5�}x�amy;��:=�x4��/����@ub�}i���V�m{��.��'���G��&�Q���Q�<�Hh�e�Ώ����������0rpz����A�v+�M�d��14��Sʭ8ǏB�!�ۼVQ>���M���	��_ti	0�R�@o��k����C}���_�]���X#Z83{����:�����og&��dx��Ma�t�k��#lGRb�1�p��Ʒ�u�2����J/tSҧgi�&e�Gpz=�[�Л%���*�NK�I�n�O���Y?u�^-��j~����3��e���3�L�^�0g�g������r�2�$<���xbHM� �p#]E�a'G�@0������0��:����"�����D����rk{�K���R�nVH�Dפ6�U��P*p���c�N��MY�$OSr�����>Tر6��2�\�y?��Hw�^�ws��_�f����"�hb_�<p�b�t��a2�u wVD*��}}�����jS��N�-V�3��&�$W�m$�ON0�mK'�;TH��Z�4R��E��vN�0�����&k�����Xa	��vm>fg�mQ� S��Y����ܪL�M�n­RȲ<��IrE�4db�T.Θ��d�U�����v׊�4T!+��2l�*��tw�$H��]X
5���(�mmM/v��`�Wv�1s�F�[E�Z���pㅳ2|�}���C���N��(Ѐ<?�����^Ll�-S�i�Z���p�O �@I.����g���ȃ�2�|�#"�{��:����X�pK����S�as��xY���$�Wl�F��f�*3Ҿ�����ԬF�3̑��fP���2��~d����n� ��Ak�~5}�����/N���X<�~ '��+���x�ߏMv�:����G�7�t����VS_Y���)�Ӹ�e�2s'ӧDze=�����˺�Td���s^�I��璝46�H��\���)��a�}Ve�IOj^N�`PT���n�ʃ۵����ýu���'�8.�w�a�p���\��n�/�7鸅��fv�˭�(�渞 *;����8M��;����v��c5T{��|���D�;��X��)|�*-T'��l%�Q6�a�2���.��=F?7M܅��ǯ�GӜ0���<�:m��w�ӟ�/r8_w�5�w֤+uB�l��{ޤdk>=�ey��vd��M`�������eB�4����|��sd'�\X���V�Ó�к�ǪN��P3��~F�y��lqc1�������6��K�XN�p�����[*��@��iJd��f�y��%�] ��ؠ�T��aK�!jۯ�D7V*d��7������k�-�ӱ׽�$]7�,���v���-H8�-$}���A���ƗX�p}�2��Tpt���s'2���8(��g�\�k/�;_�ȷ�~�=	r
6��!��~�c7��X�4�G��	GU�X!��q5<�f��dM5����oC���Q^̂O��M���Cxo� R]��.�ٻ;��4�D,�2��ܯy�YQ2-����aҮ�O��W<�a�F�F�%��Ύ���$�6��t�>�j؀���e���'�$,߾���1�T���Q��Ł�gz��/��
���(��P�*"r��rA��:L�秛���C��t�t��7d'R]�]<I���W�1&���_�c<�O���o�=����m�=E���c���'�P�k�?CϕY��|��˺�S�J���W)�*G��okn%,���ڣr��~Z��5W0��_���,��9W�����/�j�ip�L?��y�SΚ�g�
P^��%��T[�y\�(M>;�Ur��Bq�>_��b�x ��n��S�
��$��m+k��3���j�^�ď�GR�q��p�^nrz:p�6���2.a6�w�rmiR�e�����)���SA+I��G����d�vQT>��w��V�l>R\s��`OG^��3��l�����cc��!���`�Ho{3)�quӥ_�8���=�x.�@s�<%���'>��f�߱���FtGi�)�3��ޣ\�����L�T`�TF���ڸ��k�tE#�L9?!�yh�V�����ĔI:C96)�d��)��}���|��Y<$�:�21Hq�\ָڀ`&c�,�y��f��)ʤ�p���1(L�	/�)�?�]=���bh���P̗�=���:a�n2�L;�����xn(��V�Hbd:w��uO�E�ȝy�M��6�,N�nDD��f�s#x�Hh�%k����S:��~�c���jz[���V�	�̕��� �h���;��]��@充,>�2��Q�Ϯ(���j��T:�Ŕ�Ⱦzx��k���ue���Q*>ц��j����v�b=@i��qo��A�N��9s�xO)~�]m㛲�0��@��}���l1̊C	�y##�ɀl.��C�,_?�+� �����d�w�Ǔ
�b�Nn>�3b��=���o���9�=�%����H$�A#��R�d���R��1�Z����J�F�0�e��I{<�S�@��t{��J��NW�˼��<2��ɼOJ"c#Rr@~B@̐,��P�S�/�4$v���ó�����o]
��<���W��/.8'Ș��
�C��/'o���y}@!�V��Q<�o�E����s�U�S�Q/�ٸ�59^������Ջg��ٵ8� �鍃Z6���(��1�N*J���w�BE�u�Cc	��*��+_q]�f&`7}��d���F��c9~eh>��M@T�����}I7�g�ՄH="��0�=���ߝg�gz�#�(~q��E�(�RP+�X��'x�Zv��GLc�J�fZg���XO�K_����cYY��O�L��$[�Z�)�H��4�T���Y�	��/�5d8�ǘ��.冷z�n��PB�2y����p�M2D���T_�&�	u&��_ Ϫb� �����K!��7|]�*�����\�lj &<b�ǰN�l���X!֠�y�o��*�zJ�O0A�@��E��E�����)�J��F��8�fj����[��T,���R�c��>�����+"����4FVF�dk $�J�����@7y���B��jez#�������k��T/8��+$P%$X��<Fٹf~ho�ЂE�R��;� ���{WjC���5�bA��V[D�W�C�=���ؒ��q�;b�d�C�p-��B\_����j�qqA yv�ex�6'���3|����K��Q*���K�eכ��9����)餶GZp�>OOLr�3<���`�>���V�xv�������~'O��`��FH&���hB���HA_ ��$}D�[h���\+�(y����4�a�$If���!zV��p�]�xXQ�&�j�����_�2/�-Hu��!�21�����3:�q�Jle`�f����,@�I�1jN���v%0��p���{�/?��Z�2x�~.y�o"��9 ���] 4�)q�6��:)|�&+��[��С�pՆJ�$W�\�Z�D`��5����<��,�x����/�U��qC������Gy�{h��_�`��a-[�\�*�3�����)��0�+�y&P���%K ��x��Z~Q;�L�	C���%{��|��c�~ޓ�6ոQv��޸W�1� y*h=�q���@ �C�  I|li�����:2Y�@��i̔L.�|H�{q�%��-����"'MD�V����Ke���!
O;��"�9�a�<�3&cj�83%T#eq�r�}�T�k�>��Z�1��"T�ٞ&�Ŝ�-�\~S�fyԅ��[�(C�h��x�~�}D��H9����j�GA����i.j�{A�t}�]�k���F���Ois�]�r\��<���769�n[z��Z*d��#�4�f|hw�ݕ�d��)$��9h���4l@�/~� �m"��f�RY0������xr��=�(X��xp�V�w���.F#�Ӕ����O�=��m����b/�D;el;���_v,n�y��?��{(�6o*(�T��`��@ż}Spiĭ16���wi�Z� ���k��QW�Z�����ۚ\h�<	�����-4��&�!��$��筒N�k�3�O�|Cb	��9L�fB�8�D'lN��,�|��+��'�%�U���n��{�!����3c�3-� j�F|#��=�k��]"���k˰_��v��ʈ�s_�/���I4.�OO�&ĔKKR�M�LCt$�KŐ���Р9��;��3S3S�.Ӱ��R�e��Pt�ܺ,��t��4<�I�b�A����&T�a�7�ԞL@�z�_�N�[b�c	�vj���7���9��xtt�
�Gx��n�N�2�F��HzT3o]�E��X��6 ��W�~8yQ#�̒N&����+Q�� 	%���>����泿.�d��@\��'f��8+��mQ��2�2�\f=q�0�X��a߰\�'zIhc�]��^Y���ٮ�]����:eyB��jgZ�
��C�W� V��mn�(#m9m���a�?y�7�#�#��/�u�r�j�0ۃ�d�����nmWG��A�e|��g�D�/���C@[��S���>�Ñ�!�V�>����t�[qy�8�]���G��e�x$����k������=x�Ǥ^ԓ�9uΠ-W���/}�Jw������Uиs�gYBv��!���^��z���Of
[M"��M7�MR��ݬ��p�-��Ag�P��L��\�����T�eR �:O�����nߙ�`��u�lV��2�Pym��f�VP����-H�S-�&)z�Us�����
r�ZG˛Y�5�SO���+�3��h���՝��_�7�[�����pvy�k�l��n��^ô�
��5)�`ة�o�p�ӛB��t��!'���C؁Jn��6Mv!@;'0$�zqc��DY��o[Vm*ys�ʹ�UO�u.�6A;i��!�9+Ud�V\�d��V��6(��v�T ��?V�3��%�9.7/I�/(rV�&��sh�%��^'O4��7�8�Bf#�Ѷ��k�qp�.� I%���ϔ��:t$5PgeV��x�ɾ�����������Yrg�:����;k���X�=���Q*KGa>�q[�]��1�E��g 8ѡQ�y��TM^�ܰ����`c�3m/�ܝ�T�7�����Z�O��?"	D�\��s������X����2v/�������;ی#y�V`ne���I�P!M�����p�:9(��]	�m6ܕ�u5��4bQړ�*i�k��q��"{�����_Sc�،��2Xj�1`� @���W+͎��8)�%����S0����O`�iik�&�HB���HB��(貫����Ǒ� FE6ys�E�|�#����C,!-|��&��%s۹��*Hd��"�c�o���M�
�բ�~u̩yrW�QQΦ�{ޢʹ"W:�i`M�;Y��xV.��i����am&���\�i���VI�<[��8����3UN�M��p�A\�(�*� \�ˊ#m8&D/ t�g*���
�[�9_�����F^ֻ�Q˵��0'o�$��s=�)�)H�ȕ�Q��3b4�_��}z8Q�}8q��\���(�6�@���]�:A3��K�y�
Vb����T,�[�DP�J%f>��e�8�E��i�H�ȵw��[c�t|��K��J�~Y�_<{�#�d2�vك�Uß�Qƽq�+έ����D ������P_e��BC�?ϫ߹s`�d�D=~��#�orW��G�3�&\!w�Á�{��<����s�s� �z�@��;c7�l9�o�M���1'���0����I�Z�vr�l�(�x$ �j�5���)�kaJ� qr��m��v*:��>�J�T'7���owA����P�O$��� �(�4�d^\o�'s��d�a9ˣ;��X^�l	
��k%��S�¶�)j�#�냁#4�<���Y��ïfme�
�yۏ��R� ���"���nώ������E �J"�~A���p*v�%�f"�[Ts�8��0Ӧ���F	[ʳV�+�!Y�~]�@̆�"��㹅�#�WeXP�iƙ� �#k�d�\`�c�Y���1�n��v!L�^���+�Yd<�����0������(�X�'�.E�-Z�A��K�~�(S���Z��$�Z��g�&yF��䀦�p*��\����� �������
���WRff"_���vq^���	����ߤ=<���J)W��(H"�o�x�q�}Ќ�E��%A��[�Iz4r�
�^U��P辪���z�����b�e��Ah���	*�ʝE�����E�,�>%�iD�cv��;w����cVv�mI%�M?�>�:If�S�9Ft����u�h6D}��Ǩ��i��t����*|��������㓔�ѓ7���
>���Z�,��o�`rҗK)���Gx�5�'	��T4�M4�9%p���Hݭ~R���������ŦjD��:b�����}�2n`�_���=q,[��P�O?ί�"�`Lڑ��@�y���Z���g;H>IK�}i>�zE��j�t��=*H�;�*�ϫ�9û���b��9��8��#,@Ʀ����ya�a�Y/�c�.�\UէșP���G0�"{ �� /�0 �Pۛ��/TCt���JƬc7
M�J����ۜV~�'2WF�֫�HZ^r��j�g#	�O^
O�m�f�{'6o*�{p(��;�"�)����	S?3b85u�Q4'�\�,���?�;�lBn��(V��X:F+��tf.K3
�}���a�w�l;�P��D��p�sIpo�X�s3f���G��<Z<􅳒��-���,������?�"��it�5)E+!;ң�����w�����W��M,f�]
0��3*S�ʝ�����"-��z����^�b�;��"WZ:xa�NN�q1!�W�W�� �b�PޫT��d�.��2���;�p�?eP �����<@�
<���AI�� ���V�و�n&� ��(��t�Ӟs���Y�cѹ'֓��^p�M"jy�G� 6<��<DR�$VR�BL��~��s��c�5�m(ψr�)i߹�[�bS�"46�E�p-���l��h���B
���uE�ȸdw��Of|sVi6�ή-АA�0S����h/���)�O$=:e	"@;G��^*zGvȹa�,���ޢ������BUC7?���N��D-���1�o�É�m��Ǥ,����e�e�o��,Ly�mN8_�2Pj�	����!��|A۳���T2vbJ��rz�|��(����'2vg��D,TL�79p+i��zxT�p�@�2�-�|�%�a�Ɖ��C���2�����3����5�d�߸�	���d�:g�"����V���i�m��s�5�x����:�wu���+W��� �;�d�2�i����t#{A�]�F�T�^�2y�1o8&``��À;��>�h�����|tN���#�S�#����[�3˾������﮸}��O�xA+���=��u�� �<�C��Os��4�{"��m�V��U��eb�E����D�xJ��]jϘ*7�%c9q�聦-���� 3��g�-���KW�Α�5�����ֳkYU��.��Y�h�2'���C���s��WQg�l���cg��	ɇ�u�+��
�0����B�Bi��<6$��e^�e����x�K�oY9�~�5+���a7b�Y2���@�0��8����_����\M�d_g�VK�Q��3�ۀ��OɪРh�K�?h����F������(�eB1���ܷQ�$_�T$���4)S	�"�k�����=HH��\�9�~�m{h�?Z����@胦FĲF����X6#�OJ=��hAp�_O�!�s=�m�D4]zV�/���;�ُ��^�,��:��"�Ҽ`�:�V�����]�hb��O��{�Scʿ�p����%��|̎�Y1܅�TB���ƫ�BqGsCm�w
���F`�S�L�.���e�ᶷ�y�̇y�p|�*S@ª��X��SiVL�
n��!j<��r����1a��`�ҍn�]�ud���k�%_��z���gF�!Tj�Nv�!�A)I%tz�2�24��s�qP�`C��M�$OM�40 #ݻS濽F�Mj��)�ә�J\udҹ��*K�ċ}�b.C�9-��E�t{R�])�M���t�k�J�[9[{uS'�n�W�`��+�8�����}��,�a	�O�hBֱ�$AbV�P��ϮM�:uQ��� Xf��#cD<�H�i@�,�AW�R�f�H��t&���κ�]�EK���[�Y����3�k�=����@9�[^Ax���� ���p�$2'4m��P���\(G��g�T6��U?���R��ǥ9��􁱇h^��ʎ��%�6V��P+e>���Zæ&@zΉ������I]�ϒ��I�H1g��upQ�S��x`�l�BpAR����C���/� �<0�޾����68��!%YM����~���P�B�c����dC^��^1�B[3���ey>�������bF��]�����V_4�	?$�⿞���l�ﰠ�'�2�eU@F�ӼU4�O/��N-b�H@>��%��{�[��'�z�Θ�
y��خ bK_�G&�ȃ������*�f��J�JFQf�w<h����������b�s殼�`� Tk���j��`s.Ŏ��]��;�g̴83��m�+�by̕:���fs��$v�՞;/�h_�$u�#0)��l�E;���$xy�5�a@^"�z����J���<BϾ�6pM�C/��>�m'�З��b���ZO��j-+�|	_����ɖ����������glL��<"az�"VQH�`&n���F����e��T*�/Qbf�xFc/���e��˘@��S�����%tNF0]��j�G�� -GK�Z�lʍ�CNR��y��(����*�#��m���
v[�Y�^��BmԢ��'����[y��eG/b����������Oe`��'a���b���l�z9<mz�^;�L���D�ii�n9X����Ķ��QW��T��f.N��r����i��]*\���M�|�*>u���z���{�W���׫ك�����9��3}kҷ*����Fr݃_�q�2
�2�̀�x8 ��k=���6��&,��S�T��+w�/�`B�"/ăw�W�d~'V��|�pvqѦ���a�UeU4����/)���jh�X�@�Tl��W�>eǡ�֨ ��êÇe�� $�Y�����/�v8�����4Hë�(�LA�E�9��}�%RuLc���X���4�Ѧ�7�+����L54=�p���yfDO4�1�&b"<�y���bܚ�W�;�Ƣ��sֵϵ�a�@9�{[��q�8�T��諛����t�İ"h�F���O�0"�s����%��ңG���P^��@a[R)t��Τ+��������_�('H`��NK#+Qw��R��b%��4�� 0n��w�0��c5��;j�N�?8�p��X�^%m�o�ꈿ�2svgc�%�q�Xn�j�piv`��r���BW'��_�)�~�ܥA�'��-���i/9%�_���&Zl�"�I��ҽ��z���^�W]�A7���OnB��UE3r H�,I�v ��L)�p��IP̪�8G٨+�0��a���@�2��njX���B6�����=t݇��S��}\�8�0��˾ڳ�+��I`�B����N�R�y#X�2�5}zT��d�_[&�Ur���:��n�	:��t����vQ߆����ā��_�	�E��ݕ�u�v�T�H俻
���Ǽ�c �t 4&���G���wge�V��E~��1����G�$�������Z;����S.��f�^��-�h�u�D8+5��nͥ��5N�h>Ç$����T�͔�;��f�	�i|��]uq�͔+�cv]8{}[M�^*RkTx�Ӕ��	X�6�4�o�-|7I�+�rC#�LR
�
�-��K8�1����&��a��3��$i�������3dŖ�{�V�A�Oeg��r$��ϔ���_0'�m?n������G�T�5�"����Q�:�x�zƢ.�r&l[nI�x�����+�i˭c_t���f�g�*\��|�"�P�m�W����G;�E}����%��?���
hnT�QycI�w|�)�����K#� �YJ���hqb��v�ٔ�hm��ݻfը�ͼVW����e�å��Asoe�MAoVc2t�xB�4\z���^�p���]��	T�J+=�������P57k K�o@�J�ʐ-��q�J{�Ec��t�9�;����&i&�d�#��$gz6�]|��B ��n��9��pQRRt�8[:3p�4���A���X��8���N7�RX浦��wF�S� $��o~~l���K ���(���O��"�����S�N��*	o�ҍc��������XUo6s�s����r?�	|�Q�`�a*E�j
�YmS@�'&�<�Q���!�1K�2;��T���� �Z�gL��I�& �nY�x,�iF�-V��z�X	T��BGV�ivEٳ�ȃ�%w�Pk�ٓX�Rʊ�x
#�6adFGaD_5�����+�6��G��i�!p��ޜ�擽���ap���R���WRSS�!4��ܼ&�0�du2��-�L罵�/s]���8�[V.4S �,�U�+����q�k.Zr�U��z��/ MrV]�Ҵ"�)P�c��������F�qޓ�|�h��J�l��.�[GO�T�r���+����W�z�i�.�o�Ӑpc�M�,�\�,;�Xq��s�|��]v��%�c�зu�V�%"�*N*��6�6������y�I�H'F�G���"{��P�G��e��#*���7P	��̀7C����Tm�C��}����q�އ�a@g'-ze���Xti���*s"�;*	���0���8��o|l����6E?MhF�hf)������Y�Ͽ�eWCۣ�����d
9�A��&��F�s�h�2�`��pۂ(�S��������_�#��U]S�#��6{/����:�������[���ix������r�ZV+��������,��q�q��xK����&@�!��۠�-�_N�9�j����ve���sh
�����M�P݊5�*���q�$��K�rj�r	3N��p�����"ϐd6�Ɠŗ��g��Y��-ı1��'������r!dT�Sr�G�͛����JՔO�S<Ȍ%">P�R�[��y8p�ޚ5���@�*�	�>�V��:3y��̿�BSO�ǚ.{�ጞ�N�#��c���"��ku�;��a�ѓ��N�9��w��,cjp�jX�]�@�t��)7���`�B���!����,3���p
��w�%g_��E��[ge�(�_Ȉ����3�Q-�-�5|�mȵ�nڊ�?y��`�fQ���5ǥ��p�����}�T��dJ�Y�b�
)�>ȟ�q);D�A�;˪��Qq���e�:z���Q�<�9i����寯�z�Fi��|	U���N�>Z�%\D!}�f�Xd�iݿd%�i����k&X�����zӉ��m�����4n1�4���m
�E,2`x�'�)���vU'H�ܦ�C	�?Ԃ����v�T����������ѭԇ��MaO�A~`�%��ݭs��3��>�wẽs U->K�_}��v��͇F��Ka�G�����-N= u��R�2L�$!c�RX0��;���<�	U21M����
��"��ܿ'�����&w+��[�%I^Z��P�^e��Uq��dҩ����AS��fs���b�$+��(�O
5p�������d���ʚ=���=�|Ni[Nk���xjjR	�XS}���PbW8m�J��`�\�D�5��E��3Z����2���1�j��*��*�ĳ7�v�ڷ�Z.�ȉ.�Ü���A��{�5�	�TL,v���Fre��w��s.��v֛�?m����1x��b�p����N�q�	�rڙ�w������[��;=���@t$��aE��&�����S'6N�O�^����Ǡ��Ե베�&_���y�+�	�fWɒ:jG�¤m��n�ǹ�AF�$�d�˫%�`RX��,e�]4�0P�D��~ݢ�AiK�����l�1�|�	f���[��2�U*^�����L�N�:��-p����jhYH{��ѱD�w<��Eu�Ē�~�W�n}^�n�3�#yU�l��iyF�4"��C�[ Z�����8r��z#%��w^ �\k҉�W�n��#���*d�m�mѿ���2�~���l/]�l���05v��_w��&��+B+�I����6W�擅q)�����/��N
}��\)?B���5�ɑs�|�Ilj5.�rŊ�^�c���k�A:�:�K���# n����|�:�d}���K��_{ ��9W`��M���w��¬�ep(\���dFN���}d���u�_��,c�}8I}]�I�Z
�EPFv�ș}10�z	��~��B9;��>	[��Z3�$���3�-/^ ��&��C�}���+��A�/�ެ'?6�Q������몬,�2T���>Dsⅼ�sk:&3U�\tYm����j��ge��$y��Ru�E���>��Ve��֘���im³(�P���l�� '+�"Ц���7</�v��-m8����_�#rH�e�|g����Ӟ:+ʋ�����ܲ";�/M��8�m��C~l���!����C�I͉�m���U0���M���U҂AB��Wӊ�`��}����.�����`Ap��R�S�d�	�.��:����U�A��My��igdvҎ����BкSg�9��=u�rN���NdF�n��P��Ko��☟�#`��]�c���q�@��4/����Y�k���y���ba������D��jZ�9͐;x�I���?�F0��ܶ�{��>4J���`<��`�9�9f$�61�E��f�E)>=������K����Ȃ
V�J��cE�����@�O'3AiPٲ�^G��תX��;�:��0���������,��`07�Q2�S��>[f[h��Y�5G�ish���־��G��JG-�3�͎���Vncb�ɕ�T�jZ���0�߼8�ūD\5'dm��'�Qהg���1�tvܗBÁ���qk�8�1�$�|�e�G�d�n�~�]Z��ؕE�XK� Cn�#/�Z��b{� ��~��Jh,�B$R#K#{B�D!�	�YL���Q8NC�:Dv�\~��@�nf.=j+�
���'�����5�J�$�Hq������1&�La)�766�]�X�u�YYt�(�Ҷ�$~�ϒJ��3�G?�3�#E�Vn��.���B2�M���D̡'�	�l�J��0݆ <J�5^��(3"2��l60d�rq��g��K���f�H �po�����;׈��F�n�r�/�D�����M�y�O9vjN$t���������m:�3>౎��ŝ!����+�o�V��m�
{��ȅ��:�_�8e�!�P�}������Žj9�f�sE�T���9f�G��6�E��9P�ρ�}�?>���C�a�%lt�i���,ЁkeKِ��O$;)���p��3���t&P�\B\4m<��!�Tb
� ����!,� cB��9R���F�r������U�m�5�>�h��ؓ�8k�q���h�q+�~�eu܍���ƔAhu�F*�e89���g��I�,e�&ԙ;��>���ٴ#�U>p�d����vM:9��W��c*D?���u�%��q`	�ܿ|��v�X�&�=��ޔ:c�Գ��7���݂��D*�V�\D﷊�é��J��rT.�p8:�����N�C�87H-_�!�9�(\�&}�/ʱ�R@|
��%T���l�s�#���F�I漯T��oX��w�8��;)�E'��c���$��N*�>�Px������b��;�\��eִݦ��x+�$j���
����<�%l.���/)b飞�rZv�
�F�U=,	kTK�I�z���p{u�@*���:��!��+���C~i2�]H��T�5.�_9F�������Ap$�::���qv��/�
]�N�b3ܰx1�)���랤���~�!��b+���-XM]w+�~X�f�	�*)�v����UtPZD���OۼI�\Z�tss]�)iV2���!q����f�N���( n���x�h$����6�������j�ki��|mŇ� �����uݗ�`�Sx�?�����O�Y�����X$�����w�Д����n�+�\�jmmy���
>�N������b���uSޘ�|1��0ҨCL�{%k��5c�:Z�ٔ�D},9n�\!7���9�?D��re�n�y=&�b쾹Y�i�.L���d$����f�"�Gש�tA-�ş���YY���ñ5��v^�b?�s�ɐ"��B��f,�t�G�ǚ�Y��X�@C�bJ�d���o��j TR]� �~xx�QaK�1*��^��U��V2���cj��A�T]A��$�Y��ɖ$�}�D�;����F��tЦ�u�M������w�"I��V���"�PK��t`�T�@��<MR����㷎��T�3������,�X��`�,x.J������V��,B��G0����\� ��z���<�c6�Ni"�1+l%@�d���1V_%܏�}t̘��d6���;W���
ï�!�}�ʌ�c#x摔^������A�ix@ɓ)h�E&x���+[İ��������9)��Q��f�vo���2I��L�^��9��7�����Xѭ���y+!x��*��9eFPp���-.�y̗���Xp�>���Nc���&BT��� ԁOђ#^�D�4_���McH�6J��]��~�}e;�?Ψ=�k�4'T�L��4�����+A��P�+�Vt�R�k`s���<�DF.��&��j}*�Ð+�`��@R���5��� Xк�F��P��a�1������&K�Ct+ƃq4�Џe? ���$�P�=���W�P{��o{�r20�Oȳ�ZH [�5��cn��Š}��CP��$z�'� �'H��=*iR5�&9c���@����;����W�n괗&�jw�X@3��S�za�Oj�z8ƾ�>������]f��"a�sGE��.dA!y{e�(�ʻ*����%�ƛM�a7���R	���<wl��L�Ӵ|@Q߸�y*�6V��V�g�I�v'P���p{�G��q��v�&ć�������,��9�л	{�c��kq�7~�?�\�_uRe�}�;�I�%�"e���(�;�+�{cEC�09u��L����5-b5���as��4�g�K,V� ڳ;;��߃��V,�����Ɍ?*�q�(�Lk��#�1R�l(���I���$�Ȇ�D�Jܓ�F�����w?(���#P��'*�!�ڥ����X�JK\r���c���@u�������2��[��l��:�z����%�;����!�v�܊�����M�Oĭ8��������h2��4}2@�xR��7�ʴ̆M-w���Ƽ��@�I��vޘ��L2c d�+�ӷj"ZE'��R�R��A�q@(9��k��O*"���2���Z�6)2���AK�'19]?��T�ƴ̝���C�S�<^��I����~�4�y#˻�/�R��7��&[J���z���.��ε�eh&ر^X*<�/�I����u�����G�3|�D�/
���a2]h�5_w�I;O���=[���?��TtT!7�6��M���f	�N8"������Xo�D�}�k�#����JA��c4�7��6;O��|�M�_�#�� P\+�E7Q�O��*?�GӺ��Ξ��J^�h��~�����n�= :8��2��S�%+�^ͣ�yx��`���
���ϯ�kb��l$��5�r����1��Ʋ��9��Z� B��p������釬�#�ȇ�o��h�׿��!>�򥺅i(�ql�f9Ad�r²K�Ԕ3~ �lU�FX�g581��oi�/�e