-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MeLimBkn21WekhLJ9XcwM+trrwsuWFNksGo1pqmTu36jFfK6chBMSVC6P9SYn4IG+c7Tnd8APd43
5I+UffkCtL6f3YkzkiD75WcovifkxlRuOacpe674c3w5FcX6r6pRItq0eha2/8BaEXjiyzI0KB6N
NijCZ4K/wJOZNDEAdskC0OGDy9XYOBQLaPKqJ2oOfqAQNXyGc784mqspUXp9TG/7yYf8/hIF2bRi
/dCxnmlmvQuIqP3wnN+j+wrMXryXM1mhSY8SESVqidTO+3fKAb/uxdfpoBvLrMNc25kjI2zl6P4Y
Q0Ky+Mtz4BzEekNF0dv3+gig8nwTdki4aADdBQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8064)
`protect data_block
OxRf3aPKWP89EykcWpb3R4psL9roy+TWCDQp/aha6/etu7UpRCtJnMrewDR7L206qyikjlcOn8kT
E2ReleH19SbaRzS7fjmA9uWJx9J2xLhjRACU9rlWp550HyW5O1rPtOx6xtjZkRkLcbyPKQseyODK
1tkhGF2rYtJ6j728p3z7+S5jfT1EVMC4jEE3gqflhRVn11J0K48oKF3aSpbSKlrDamnZPveVrTyp
JeC+lGFqxETFRSiNKuG8kNJGzcVrsCro/8e4QHQHv7NjSJD3CDsKXi9b0ysGsX5JmUE1yjea10Da
8vw1+Et16b0yrjrt3WyEWRcBsmYMX7ND5ipUlbNHUHpJI9FWIYfgMAKpEX47ZGpvp1ZXGq498Op0
HSZNTc2QutrR6t9Q4aa7tuNt75BkjT4zIPGf+FsETRYWJIHxZIJ/JJvcEhoajIZphLaST5VL7lAg
fCzz32Nt/p0rE+nZ5GAE6Xy5z93GP9EuRFv1y1jWEymrdWLlD5+J9CnUtVVfBokwou6vkd9U67kn
nDxTVhlA73d2Vw0HMiNRFD4LbEkw1nycbVw5kUrOXRv7rpZ6jJ78OYsjjFQIdnCNVxX5sqeU622o
YXk9HJQyoU7cEKXrOaFh7Twel+Fmw8cTbiaYMJIBztnDnt16DZg8jdTibDcBJ6AcS5rsEGrdnp/h
wRV0qXLKulAXfG7+5HSEALhulp479FnsT/Yj/LLyJHVudc1hTZb4XKHZKX2xJK0TH1HLvKurJVGR
eK5OWeqspG84X0rCyXhMHAaNumgxQ1u0Clg8IhDzjGzkdlVctWnPK2WrEY0d/vbX+Ckb5kKT2odq
fblwnqFLVTSvs34PmO4SUHGo1sAz9UCLHO2RDGqTJ30mCBR7TcwcNtSbIy6C7z79zknzvMSwM0tS
6u0XE3fF7FkLOAoyXvydlVSZN5zYUrErZi409wD/T0lzcQerS4w69IPFDABrc6q+HdIRAECgz6x4
ZI7+X03MZeZKN2MwORvi+wTALMgN0+nCzCdTPikvyZ2H4c94rx6pnpHE/9HZkJl6b/mQsqNX5R9l
MIEhM+lQXrQv8f1IsA6YhbEugqUnSPQGWvlNHMBcBjHr3bfLV8X4CO6YgcXuFLmaPcz2uGrKjfFV
S/8r0Vhsuym3NMZgK2XIDSIKttihRCP5s6AHyEJYZrMIvdIjcQHBLVuZnUwHJE7WSb4cxpZO9K/l
S/BBeDWv0vJPzYDPwKkVYfMDSzIQ/7RoXeogRlcx7x9WNfO0levWgL8FTfpUgEgnjQU4GoXb2osR
Veh5LNE/uYb9e5xGjguMUz7SOlpsDAGy6xTSCsjCweGk4isnYv2dt6OZyC6MtB3Yt7GlQM5V91TL
GgoeSrgtPMnaVaj8UjM8iobPkwbPYBM/dxC37GKLziSxff6WnHu8tZC3e13HmTv3mAqv1ZHvHkuf
/kHEkD+xSt7EsSHo0bLbLSfnPB/8IXaHWXVh+IiQrI2JzPgOgE6oSTTPEXZB1tUdlbW3qTxJeS+k
7UqrgkzJnH/6UD3IfV01FbO7hPagMTSNdZdpZZ4560/TS9TFBGg33LUg2CxCXbYt/yJBvWDObt9p
i1Xik6SJjQIgjgldNzgZuvd4tYQb6VyuXDs1EBQtED6e2cs4KadXgDOLZDMvkD2uTCzes3+X0Gvm
RA7erkAUo831XqfQ8n6FPJynSYU9qjv99sIoIv9mdOtFJeChwoooQt4ydwA+akRqllnHBesuKjqF
YpVyyaHaZnEQ0GNyBc6ga/lcLq2haENe516grxA7NEu4ryIU8qZy0QQ3BUEq4DkQeQlNlMhWneIw
8Zc9ztvmFlNtV9ViPT3VPk9bxefMBV7OLERNUNCjcj/AqoBt13BdfpKxY9sb7smHnkBlQ+/Q65Xs
8g6AUdvbQcQmHXKHf5jZVHk0KmxvvbjVlHahBQ5MTe5NQs5P8adpBucbLjqxOqEk7+DMV8R5SbAK
DxeuWLISO+CC58uLqqpJMrox3uoyCL/uqF9JkD2hbFoTKq1SvTiC4cRgO0f3mdc3kxWKRIHybrnF
WiPwVB5KOjeVikLM8Jgvq/lndXax6O5kh2OVh9tNeXDOzepQ6RNRbB8c40s+1SKNxpKckzUffeL1
MnZVcc3U0Mo8fFOTX9XiAhqOsijfoiyU23YJeWPjpWa8oXCVplLSL0izrfsAWSi78EVJxW98bp3Z
hspjkKG4zG9xDZsFB5k+KzEtKjxPEx5OMpF5GBRlpO6+UxaYJ96e6xxHG8sX86VFGIJThaMi6N5U
0PX6oX66OTAkNtMO6kycCgiZ8K5HeZ5nRmyd9gshm03xDWxge96wnfC1xI59bfq0pCaivT8jghJT
E55MeitTRNlbwRJvah8gSuRWDyd0g7Z/5789d8YERx7tWzAa7Fub6GcbKPofSGzEdxALG9ppm3x/
G5MU53K+4kthitHbUdFxHlIh4Qk3O4iCdIhUO47aGa28bmY1dtTX2WOAFjhC0HJrZCXinVhVUwrr
rLQ0Ss7dxhHDGhS8ipKIw1AkmJMsJKqnrXgGmnzmHx5kBmES7vpH0X0uPToTuo9n3YeqIalu4o44
nP/itmdfC+lT8xl1Gi8jO0+cYN300zY9lzjQli1c8b1EjkrD44tGD1VhDbIvmLWBndxYyyzzXWmR
8Rul4gTYQzPpbdec7u1IObj9EU70H3n3GH85oVlYNt1oDsDVqNB5mRO34QnZWsiVHl49rH6SiyfM
2ksb7eUB0FXhHsrbDHvMFAES623pqZ80Mg9I+AUftJ7VAmtFulF9La/q1hSFWVh87KPfx4cVkia+
yibgczpg11OXedkZJmPY59gwDLaSaGed29Cbvx1R1RwwptnJrAhOWc9jlvMQjG49ysz4lxWd+WiT
wOKTtceIi0s4vevfyeiSd/bS+O+wU2VS4VkIBv27CQw9sEd1ZZV7M570xHUWHHdqWAiMkSm5LFGN
BBkNed5RSlktX+v1//6do7jUyAzlUINh4IC5rhDQqELLdKA2Rk4UzjTDyFbITbr/unIqBteceW0T
5PVvLuOXkGbKzLEtWr4RLBcHOn1qZ+//SSSwdmdR9J1lFkpRCdYIrStqE3nNHbi9ODeRsz4/WQ/j
SANi2gJmKpf6z2/2QkvZirFf7B7HodpR07KMpm64lb1hc6yJEdDEYXyd4+iAC/ckZBMYBvZWjAAN
fCsjVm1MM6TvigUjkPhMb8PyCO52dBNPhwN271rGfggxDtt53l4txNxZZtC8AKmvbq++ZtQqLzHr
yguVVK10i2rSqrzkqeC8x3aQyOy+AIcybeorWddimPMWYR1KUOiwXzEY5FUTZMkVXMum+7bPjmkU
A3D/yEVa3h7xl78zs6218M1yyyB12YkBCX7XNCfLRJYxPezR8n2T1B3gUwLEK9H6sM17MKM2rVHb
FbBcRUlwUEBJYDhDDsH5xZ9PhaNIUe8SUvOg31EVxkF/ZbIksO4cRDBHr82T2n9svkiVLKSmnlAP
tvxqlHEP4yY6ZswZ2QreGDAYS7LCTyTV1ylFDQwO9AG5IlWImz4SMrmA96vlCVa1jY+tEfl3ah31
SsEBMIhFq5IedoCJvPoBhxzFNCxhbGyr2GtVgUEBXdDidTFgoMO0ORoXsagI2d+HhGAW65qrKNvB
qhHKtOG1Fs5s6G0RgxTiO1OirTPaQVrbcng6Fl8l1UwoqGNH5kl2oB2cYTbYh10uURzF275c+gNi
9N0hQfny+pbW6IA2Xnm1Lzhsf6Icayc4sOvc51SH2kM98YmIEA9JbJ+Ke5JFMH5kAD/Y1/i3ZNKd
A1NXT6bmp5HTDDtroIjq8sgO/iB98swlzESUgtIU8VH7l/6gKNFfunbovxGAgnC6TWo1c2Ot/K18
ultooLrenHTrQqY2ev/PXaWMnw4dXUKkLkWdAtvx+tAmyaiZQpfCxzCq6m+Jvrkr7VJeHLKK4p9q
Ttds+7rBrfaNJgOKBhJOrUCS8Cq2+5cajeM4Y5f2IQ97Kjkz95xxuIPW/iCOZhiPt77zQBxq25xq
NwCOwpZc1C98DE1F9yiZjxZiyz/kGeHrNPZxQSvNdi/hIK214dDYFQl6rixccC4r/QGJS+rknBi5
eLxt9TsqV6x29NpK30TbNzTch9+UHFstNr1d2pz8xmMawl+JZZyd4gL0szT3xaqlqau0aUcDJnze
9/fEndqkCijY2Eu6IT7lJbsdIvNqeg+AQS3a7yUE1nhm7JfovLYv2ovvFS6jxk/ioEZ90LQvZZZQ
1DVOqhQOSjRZCf7ZZdtTFS5fjGBdegh8g2yafawG1DMe36ej6cO7oAG6htvDJanhKss/RTi7x0c5
+8mB7EfNtFnaKKY1N0gFf2Gb52lKbDsXmrgD7XA6H6qU6vlnEsffFdPR58qHRcEQrF8+h6sg//Lk
aohthxPvdEbi/Fc9N2QsFdChAKe4ePCROMFxn5a0Ie0CtWmG6xAcmVExaW6BwnQ8MkToaZPLfzJx
gubcs1emRO7snm+uflOdOzK5Qopk28ymydvlORbsLyeWha72r2rzSp1SdlTC6h4WiVCPifstKP97
Afq7OQK3WfZ4OpQEX9Uky7YrUUlLP1Hz2w+aL8x5qD9irkQnGxKJ9xRh5dX4vNmaC/1b7CNo1vxx
ezJk7JKxmRNgVz34TtG3GKBWquz2ME7NxtoQ9xSFmAhSOvhld6P8hBX4KHcr2XRmybiHiOcCByX2
I3ek1hjHwJ/eEvedOOyj359KImqfUp54m+EPsz4vD6B+zW5ZRqyckdk7C9c5eN8Jmqcj18Z9zkUj
15gf+YgyNJ2xo0FJCHZGwt7M5G09rDloOTVgxE6hJaA85HKWMP7uYrEJ9Z5WaD/nmnPyUwMrktrd
BHAmwhB/a811T9QlKjHz2uzXVmVTnxQgX9VJYss9J+bD5carBkhpK3xgo3yFHyeh/9dS9nyi7bvC
lGfq6B7R6i8mMqXWF/5bcVgsO83Aii8sS0ezHDoMGAzDkPbt2GIridB7URterVtY6Nw2nAJTucpe
jM6nrKEIK5TFEKLAPqdA1uPY9bY7fPGj2GX9711F+BYa1yZwOcRGsjf49MY+riA9vpjywMkhcOiu
QTdm1W7hWK4HzpZLoW/obMFJ6HsCIC6lZnu/Euct5B/zJttT+1vvhvQ2CJ2NS4iGSpFiP1b3hjKr
R5kJjl5tCBCiMk42fWp/7QhQg0DQAun8+9zGRB3NreYjocBL76Vti403HAYMoNTN0Uzw/z3ytgHj
N3m/NZqcWQ00RoWXx4BrFBo/bUZ70bihsWQEnu43R0qoEm9SEm3EbfcaNDM3c+CvZ1bV0B79fzLk
hJB7U3opp+afwQfyfya/dFoPEuxCQoFJNUHgptc2zgoa35tKX8yp5aXmxNyCyd2ZOopOUddXch3d
g/T3/XI6Eu97kIhN1JtkBrAS6l6yL+Z+C5tEsMVqDEpJlXAGoxTYYDBx8Uj8fksZvP1EKURIrjQQ
UZ1TuABoe7J4a+2nF9TKJgvScr0hYDEZXqh5/SXNrGcTR4z+PMyQGLD5fkFWK72V/+ZwsHi+QiCg
gXcmQ9j34Pj60EbrziYxjyH4YK0UBMyrSw4VvWVCKen8bP3DaX0enF3m3yYzA2QbD2iHucjy801Q
UEPvTiIb/IuvxtAl2Rj2f2tZN/Sc3HaBFW1AaMN+YShrEzlgLRWnDeQLblDtbdYP4l2zdQjq8Z9y
1+fKMRz8vRAGdldPPeiW8I5MTYMa/JYtZkBpJWfdVFGq3/TJjykXWRUez43XdD1+W6I3zkDBokHs
alLPQwO/23g4eq4RcLFKYJBLxCr3kzj/YDeGlYK/MJd9odxlr8Io7nC52FlfZ/J0LLTtflyK1bwR
HfxpLkPdIGxb4WtzRkNRhVEW7di94ejjEB+MC525tZELTaUwZmarmQLLULbjrn3xmSmex1GScUO5
VADr8FPtsBJrAnC3kZWJX8OH39EHuKlMdZsjb/nkSlLAgPi4mug9A0og4HA/ci3MQkkAN2wQErOQ
7b229b8fx5wcEMOK15Q48jGAu6YQEMWO3FOpqIM1IRhV4/sOhQT9HFi18ShjcY0G+x49OiSG8f7J
9636ZbpDX5AJ64ti6U+k7TrjpcyZeDUHDpIlN8CtWXZrJvQTsHRpG7l6IhFq8uPUJ6vDRHM90Fo3
YABSQWrcwANrWFvncUxo9w7jKbq2TXg+0F2WMCyYdSkjZRxgms+vSdEZjpOzVJNcVDnuMNnwqhFn
q39cUgFb9qOdska41E+NSbEZHJ/wtXq8gvVM3F5hAlPthUaXV4oM2fUmM8cP6qV9nPKdUJWa14Kk
qcieO2cwFz65O28N11+/mn4mZPvLIW3WZgJRVEoeXb2LEdScAkkGL0G/wINWPpyq4hMvLzKQJxXY
CjWY5H0j9izCepxnoBEE/Mcy7TQIaLDPQ24Hz44aSKCnA7IiURh78V3qn7AldklH+UUDvfGbwIKE
zNM5Z53mxL7FayU1TS0qDb0Mt5d++I6OiirWF9czxZ6bgF3tBmESGgFBnmBzu3xIyMPiCcF0esQe
ob8+UiWNjXLB6mLCjWzONnHtx0qQRl0XY7n2KLk8x89tRZy0t38GT9ocm/PAuvZXxjELvxnvMi3h
wyGs0ajTgWiGIBoEN6oMrz1p89JCby2DbF61uRtynLPLq4Y/fwVLSqcXUaeuM+VJkXjNuH7m7Fus
Y7pXYUW9+SJXlnb4eCEz0HTyv3hPwzT5exHbK/fdeLjxxUHA9BcRSKcRIAhOSZWhXL907vz26uFW
NBfLfcjN1VZrVYLZOaf9BEgHIJXVpWQBCnuowXCXgOciCZJ+ZvzbtoeApNVygnpJIqoEIgbU1wjl
0qRj3xYQQuEpMcg4qepPwQUResN0ydfWX7EegsUqF5Bc/riBtqfq5HkDWQv6kzsfUMXL2etDzgAn
DhtptdgqjKZv+CnxSAX/y5QbT4H3zqVtOEObW+ZrYvL5lCwd+uUZQ4t+bj/2FqmJDJjlMa+sDBp1
cqo2vGYqRQ0kV6GBD8IjQoq3ieEh29yFOORP85PnVJh6/TBQm4x2ZcbbgYhXI/bLeBZ2CLOrE7u4
i4j3fFPreBlAMTLPFnYx6yrjw/SGIpBJo3P4mhmvobsaCgFVfcmVUsOL1nXuECVOkvtS7N1Dn69w
hZkO8iBF1WrwAJtET/pEvaY9eLO/pkQ9nXlFre4egMqW6KuF0fIuDvb5gQ1Lo3lqJWMXGVkorS4n
kwCyca3JGvo7sf2hhTzhEdXj/b3JTsAl97BiCKlQzCQo0eKiZtr09fL9lSNQLRKOLS1bhkMPMJIj
rHENls6vWlReKUvlnP0Hmo4N6+ETkT/7ee83Jh8IuvhXEZzkXZHqz+0gxGXImEcR6fdVVEvt0TAI
COBf6loFhbo2nkyXl3N8mGimfJGAjArqeByr74l3lW8sTiKN1hB+0lyZqnkBPSMr9lCfKUOxU3v7
+qfWEV4K0Ba1UYPxWDGIW8wX9o38PDQWBWyXOIw21H0wj/w/mjzdkBxYRrWWIJ3H3UYSzotp8CGZ
+ypcQRRceQIc0zQbpxrVeDDCz/Z8Kq/eX05oFqcVcEl/9cnfB/of3RrNuSb6Fwvgt0vXFRhM8394
AukzhbzhGl7O5K9MXKAvd+U5pxO4TeBezhNmlatJiG2OT98i96yvYVcG+LEM/ct6Q+DWvdgssIVE
lk8S6F+ItlBgeIsy4O77IaD+fdiCmjHAY1ImWBfacJRq46ipVJPfoSf2I1tHloOMDJ0gQX/FJjUr
keFx1I1Nu2v6PWoOEOYFIh6o45LOk8JeJ9dZFj2G5mnPGNxNGP4C6C9naQ/2khmSRDV5wzwAHbwR
q1VJup++LhW61Rat2M6bimzOE+YLCIJnpug9gA2TM+10/ZrGbEFvBjQowKi8dB7uHxyEI1tlRooT
CJIfITEv6MJzpLabv8wJkH/+eIv9PZ9bLNgGXUYLojVbJeGJjna704EET6klku8vWPjIsVINmwKL
NqPs420n/2Al6V8zxhTehNawVFpipSnjdRzEXT2tkd65wJWXzeA7YXfSt5AwzeABpnE3X18soqD2
v/HqE2WdS5q1M+73txRUEC3ZtvVIYcGSZENdj/74pFBvKI6AcmEXowED+mS0cjjUK+BlG8/ruPxl
4ua5bxtL48GbKJ0nYUNbFokYozUxpUfazWHis8OTAn+MGL33yezZiRndEIpsE68bAicz6/HnfKSV
YSvgVSXTujyczwtCGdhtBRwEsXgpC1AVmR8Ss8N6ykpTDrPDx48uRa2AvUNyfPAKGM7J9ZexObPG
syyg4rL8BhB9REHR63ikKJtx2imgajrAPGtCAIJ1vmRTg2MGXjT3TJC16KjGL9MW3gzROfiTKjel
OBE2TrHTDN+xx+rSKE+iGpQIy4wWo8f/3OfI0N5KidUX9Nttdol7BnCm4IBrhyC7ZamhnZeVSKlN
pYaFFarPqYyf9nfftKzBKboO2eaWpvGsPdup60GiOaoqzfwPXpFTYlr1P40dkjJ26sCUDvwXBYzS
2D6dgLpYeOmvkxdvZYCVIGnGCbi1hSMhMBUH3XVFUNkRf4rctzP5JZL2952Kn6044pBDJfAw4bTK
LIbM2thkHYSP9ymdYXGaiw8oNODqMhTv7zptA+7JSB7Si+wQpULDVWac9XgWsNO+argGnnT1cViN
YdGZNZzgTU9P0JX/rmAOqu+NwsRsVXxwuirDae7lOgiVcgLGWDvGX9g4zkWkhM9mce+w10HzGrfx
JavBr6qdZlBvz1LHb0aLN+mXHhgROpUcnZEvKk/5xYewk6PbljzxvGY1XYKJ6iWvdd4qP42ZoNXy
/WGJHlwzveT8pN4jVjBfZBocD2L9WDL2qGwsIry64E620edN4VzlvUyqfytpa6a0v8iOQ7lRrZF5
qr0ay6frz5mRWOT82wgXQyA2TKUWuhe1JZV96E382Tc33t7kH805LggPaPsm3Yeaj31ScVyUHgWX
TMkHEMEWObRNM34IcIGqZqvGpx7fUg92TalS/oyJmvt92fS5eIDvpT390/cXokZeWfC06WD1mcY3
T+8O6m4uRkHrWOCae6Jc17yqop94OGY/FJ73U6xm3kTwX3iUP/tZGdsU4GU0Wl6Y5Eeam7iG/NOQ
y+ULjxxusfzoI+yHLnXPgbXZGJ8i4NwFFxlsPGLDoDAB5w4X9pA8x0tTUph7X3RAxIsKZNJAnswm
O0BMLsdWL9MLNVGW2yOUtrD1VHGezRNk+S4p0DS+gJUFEOEIi34Mdhg3tsw9qpLTdE4vM25WdZjA
mxCJTkfCdaBsb5ZGBkUTms7UHN5a7nYN4dWY8RgXQNIvfNBxPsHIr4CKAYZZCHn7zFANvQwVTT4d
f3axaooJbFnzzOI1qfyBqpeno5cDUrHKnzabktOErDHwMfpfYw8qwrHDjAKbpb+ZsVW7JQvmWEHE
tEMec1UaHjj0JbUJff51ZOor+Z84YFRYuDTKplM1GccTAP2acEwKnji5vcdtyh06nNRiC1lK41g0
9lcgv8R1xfWAxOKgxPNeOjJpt4AfPauHc6DkIYLpGO9gJjp3fZwlLpxuJEY1j0FMwVVxcwltc8ur
2NNBaU/cv3K+NAeSjiPWg+L5rszUesA/nelINHOgkDIVipvLGhh1ITH/IdwC3x2llsb7sRXdKSYo
kuSzNyVuCYnhbKQB4scPl4RilX/hZwXLIF+c7cw1meIBtz2CmIUlEfdiHBPr5rO/a+DLxaF9mky3
HJDOfyOgydB+Lv9qwRcmCzCzyhVxP/N7r+1Tgl9Rthfdl75EcBVJcyZAvkb8RavECvAsV+3Gb7C6
E5AH8R8HadVbqpcNY7VtyRBckN+A2WPK2YR43B0s2Xs2905uQWnl9oevNT2Ujrgn13w9dOOKRogr
Tc15FRjTyPhur5YMNUOK0+7W3CQN2ezgu8GzcK6iXmQgeo/QkD+e8HEDQXKDElYsA+0PCDoYRmAZ
QZkj2ACux55DLl6oSg6pX1QN2+A4PkVTNSUySv8njihfHPMzpXttsfefdSH9TVDLQjjtPfvtcfBb
OBi3H8hv0wqHCtoLD+/cEikcLTf335x/Ra7hAaSpHRc/gYyc6qLkGpoEJRnCkzOIsn81e0q4a8Vc
Nu7Os8ng1L+rb4kNKh/dB1HpmT71RjscjgF7an+Q23FMhfAtQArKribXdFeoV7FVWdCu7b+nA4UU
w7uDvIgQkRxnbyuQGbe9sxdtj8WqfHapOKcyZcMYLCS8kN3BbZdinxjgh3HQstP7cZYQAw4tb1Ef
uoEXf4UOhhYG1CD+exlgA7FsJzsWt0TBsWK+W2qcRK2yZqxvty91lZYkUH7rP3khisJ1qiqzkPV4
CKMMaIGU+/1MtAA4Wh+O3iIiUF2ukbeP1P21WBzXYQny2hQfHRxumG8TceGDhL0k2jfUAke+ZGWU
6xHZGP8dxZD5eVaZ7t+l12ncZvedujdW22K2+vFwERj/l4VC2fSsRUqncB0EwpemNCbxIBS89VXs
oFp0rcGNGDuYbxct/YwKlR/aS6gy5RnrCk8pv24QuXZxg3QTuI5bfi66pbx1WMIUGdxfkLOcmlij
0t5lYLUY2k1btYD8GGQ3OocPK1aMoC2rl/00GjP0qMB3emwIqRb+V5q7H1qslW3/xDPw8BnHpeLo
6kat/kYYhc7o6ziQrDmlsXrwMx32hixH/IZGTwQiAsXYX3sv781DMg0B/ll0QaK7D5TmT6oGMPJ8
KNb1foMGuFKHfE59GYqc6DpavVR0HftgqloW
`protect end_protected
