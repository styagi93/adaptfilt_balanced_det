// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b5Pjp2zuGeMbDpd6NT4mamjPiFN/ujT2tDxK4VhsKCVcLu+vsrf2E4ly/ii9Bz7z
n0rtNHoMEN+Em4bibYRVWQmeE3k7uw6eTLL7CzPyqHpl07TrodEivlRNAjYttltw
H9rcyhgMuH4b1oVbpf+NbziZlpFS6zssxssZ4Wym8mI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3056)
gGm5oCC7PDoItMmEdco3y2W1g2CcOQEFytXXnAJBJnsb+FSel4fTUpDaCdJ+wkSb
EW/HjgHASFzm8HtOk2IL22IItIRGtXUXmyeiuXtgeOkvU22kpnxmgz8FqNJAhwtQ
mL0UlhBq67vkv2bUOhuvjPAQGGcKhcqegTzQFyWRq7nxF826cKhZQ2NDmMXszubm
Hy6/yvICgtOGf3DDyWJPx2rZEroo1NnwZjHPury1AEofkTHvrhq8JbL0QLhpS6zO
VrVVlO2uyWtFavyV+vURcFu4DcowQWpp69nVAp+GHWyJ0IGvIMAe16c/APhcQmc9
/GOSfGuioRge0esdIdbSXiKb22MZkDJbnPJdP9qksklwQFYLAqniB7StPkNdhhtl
ixdsXACCkUM8GAakgxt8ojJ9DVxY7jkkr/N1aazy7iPD5aU5hQ31cL4eac4XRdR0
uj1TDa5/ROd6o2H1bjOCfO7t22/fFp1bae2Dp5t65VM05yFSrGJbFfPU8/BgTjj7
CtZM15+pqDr1vhboM9pAXgBcEhwsed7YvamygUZ5QJsI+KYmafYw/iywVwBbFpf5
q/exgrMIgwx0r1hMO+IYlOzblCeiw/RKmKP8//wqzwK6YAhQ39hpaLmqqdIE34NQ
8vtxLZRmvkbhsvfaapfT/DEPSeVGBrT3/PXD3FTdZdZnqH9CM5QWLJ1TMStp9F8H
MU3KHNGXU4s61IdIeuRqtUnR50tDi+9BLpkmXMW579FQJKCyXiwU+/0sHwR8DkLt
k/18ofyxMiEIuTtL0p4vW7ACruPJvjSPDP1/nZIpSvpJci+TVvchd5U17qYBVtB4
6fqDgU70ggI6C1zOX9bci75Oyq2Ia6yLvrsql5+we1fYxzAyfBbTPgBFogqnZB/k
Y9Sj4ur/PgkG6M5nd9yipe6ojuoO4GFRcSi26AFnpTtMrkvkPbYZTWHZJw/UHXwl
SouB84pFPi8AdD3VyH0DfiLzFsqD3nad1I3noY0omNiwIEpWYnpRlHjyj912oMSu
OgAxDzaDiOyNp6ApRakrIe1ZMdRIrOeAzleLhKWkaovEkmPyhva1yi+b1J6Bijns
AkD4dCmcqUD3sVyCE/bCztT/QqmKBMxr9syDmCLViasbWOqEofg5w/EA8yk6nMqG
m6Cnu7SszZgh9AXHWWweMOD7ruVnCohoXGt+JcZTI4kq4bMSMzx4hEk2xUV7cufh
TAZfj41b6nei4Jtf3JUg1z0W6grkESY+Cl4z2iSmNeIKV0FPKo3X9oRdBKdX7q1f
1AGWt6Z0QsX26iReQ/74LNhhpQKnYJYFeAXHtSUFB645BAFKdSMwJVL62K4fF1qc
rDNAcYGlBzcUaftuYw+Qw0MjOJFbC6I/bwe+Zdoqwk0uiTrcRsaFtqCt8NphDykK
KDnr/IBazU3BmAso+ma5J8jnLbP37rGD98AEOVkTg1DfTqLD1Ut1O22vdXs/KCjx
0gqEFT+ZrR9bR54nE0MJona2SSBBGeB1GVMrVDd7Y0YoXaY+MfbNAq0pFQqKO3Y2
DdV0jN7yTdSBa2unm8atcq7ya3/j+9rnIcYmppAgHnJl3AoqrCqri4SBdRWJ0LKG
EskUq3aPBLahBkBQY52+UrnWLvL2bVoaqxO1gJA+fmlnvipgTYqsXRH1Yb71U1TJ
tABEbk4ifBR6YbRr+tN1HLtUTvDVRa5tQ268KDp2G0dzD1tuQHHkvpyxtg1Cm8Se
hrMWniHOsgMVXRg6ZYZSfBPthycLJVFpCuHQB7yqN1e8PfICwmrPc2Cu7Cdl4C+n
xqm3hG2c7oolKG9I4cEM1lLbcRefCVuERAe3eEHJlNMHbKpLv7Cy7pGfh5irx7TB
sBpmtjbfYQYoJQu6TEXxohY3UXFuin9JI3SrThf65zX9LqKY+9h2/9+tQcPM4kxW
HLeZSkXSji9W5rvHg7YpCiXVaXDMbh4AJuvfRNtTVs3MIe3fj5dqzIWFPc9TQNOt
kuoG66hxqxM0uAZSzJJyn5iMVGOOGDE/gwqjXIKzMkpB/763cVuwlH0C/iyn6Mk1
j3Eot+lusUu0A6ZZqA2cuYlZ5jUub4RyAmlvPYnML/Ym9RBc2XBOKbORTsQSU6gS
jNUdbJg29SLi2TpQRcUkgbCSHd60EFkvHYDpY8Wb+jePfdZjWrblloCk81ZQYGmv
iNfhqCVhVcUkwoK0wbGU5WUD8weA8DT3KT9pzyQiAHOZnyXEVpayNPilv4Ef0yxW
TbvK628GmXDXjOHGj44CJgzFtXfcN79saR05jdgz3pEJbrr1gs3+7pN9ew8Cm8XR
xsy0M1YuIrcWw2IR4gOjAYF4uACWtJuZ2Jbt8NiRjJG0NMIRLxexSxDwQkyn0ffS
8P+lDhynxwwJIyBtPX0tzjsgf+YETD8XDcRGl0tt6UyFuVoUwLV3wGBQqYCtNe47
kva+zx5tGclfddm8kwHaRov7GcB/nHP+L2/WXhb2rFVufZKVGeuXAqFKcDRJcu86
RsF8cx9VsFlfGc6+CztlZupnTJN4ofPZsCjUIOiDC0nYTRdlIZXWL7MWxTccQe6q
et//Pqst3EI9FIVQnXdiMDE08jVrqWdwqPWHvpJN+m2AhcXxcZ8knOuXv7l2bQNR
zitVuy9DK+u5wKqRWPI1VrzNCUlNEKDd/G5NDzs7czK+Y5rqEpZxockFn/H9fGHz
t4Vf16FeKluqW+OpWEOEVTXYMESlpPPY74hJ3gtuCFCqplRiFsY6Y/Kay22f9V85
FF0Rtl/siaYZqxU1h5B//+LE4IiZhhXhd247uzw10WGO642w7El5E8PCqcSqQE+C
HifoyhAZ5xvfdcwBW8SZiEFg34Oiycz7fELmdLDJddyygLiMpukMmRjD0zHWh11P
xB+PFjjB1N1S3bMfHtNcwY+22TGiRr7td9y/CuKscQnam6AB+bxWPbykcXE5Bzb3
Z1YD2B97KsAnhATM1qdk5WGsxQsQjGc4VWrEBnldw4xTbjMO62h1ZEnLzPjN0s94
J5wIDpA2a/QFC+an53T0nTdmVnNwnr83MIytDGvFnmCqKYRzcJvsd6AOs4khfxiD
OBe5EY5yPFs+vTgh99K57rQD1vH5bgcOs8nmIi+fea9ZRnuF6GyGRdWqEFEZcPSd
F2TW48GA4fjpRejdQxrCYYTi9tVYp1TdPe2gNmW/lehL7shbxb+YQidMKrmQ6H1t
2MIPJAoJY5x5C7R8HB+ie9n5w+dKYUO9TiV1mZ3YY5+m/iivFcYNlzMXqppELWIG
haVV3sm730wWarzJNeunSONnILcsqtTV3EKcMj2PX1AdcAEVbXY9I12YwAjNeweB
mhIgGp5dfNdOdu3t6DOrdisUfeEMg28Vrl1Gt9kgOZiPafO7BWBNv2xKcOynYkth
2unnT+tdL/jB8cprTdSLewdWk9t18rn+rY2aC9dAjuMtnlOrFbWrouDpQ9XnpUE+
27svQapLIr2rM7jFRCadD5sWX0X2e3jXkvsKqme13ekjS4f5qgLP812Y6GmTIkPa
cxOWjPRJpijiU/TkMN1VN/tBuBCpENgFJ+OrvJd/xtSTuhmjHkmWybfAdWgtoe4m
TAe2o96yb6XG5ge5tTN9ihwzCToKAy49PMG1ofQOFVGigSkCr2drOL59iozxzPTW
k6AfKqBwwwjiLh5dT8FVWtF4ZbVEIlsD3mtFpll9GdLnDHs9NovDGfJfPu4mt5qO
g+PtfShUUHB1zw6mduWUdBdQ4/4qAmvjUhaPemwmywqohylShZ1RW+CVPJn80PLc
8beoKoRqTVZPUegT0e5XFiI2XwC/O+kmEL7LyZa9yJnB6IgPOlHM6kid1vkioTF3
5kq9WjvoMHKk36Kh47nK9znN1KIT019u3miD2Shgfp2U4UUfub7IOCYuhNO7iEMJ
ki6zk/2p5fNsFrGoc+kONY1fP2xgoPzEPXE9Mf3kafhCUTyY9BTBo5fTDxIXrAKn
Ckuh+AKHJYv8virNNx6tkT8+Xap4IZMwPwuH2pDJJ649RI7jJLthA26CY0gRewvu
M/Jn/W7Bp7NJG7v0Wo3mNsKKV4LGPZrq1iEJrnHMyx0=
`pragma protect end_protected
