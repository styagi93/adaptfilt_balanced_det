��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,�H��#.z����?Ď[>.����Fa��֞0�l�x:�~���"4��,3��^�?1��3����u�\��Ҡ)} ����9���a�
��[��P�������.�I�P��b��';�b��
n�u�G���$|n�A���)"{[\CR,�J�oQ��P�iQ�|�34�k�u�Mre����p�@E��Q���Ms��/�������<r�AoL��a V%)_~�(��2L�������b��P��ނ�UI}>�<�?�ӉC�3:V�ru��
�o�R?��]$�;��+�����1R��b:����"�xzWq��/y:��c3�B�3����^s���GE&�F��0�oX�|�X$��Ή#K�g���JM��U�7D6v��>&�c7�nRg[0j�C;_6������ǅ6d��fl��`��)P�0����_���7�o��J�Q�-��C��ʤ�]�m���a2�5;��U߶��+,��].A�rU2MÖ�+����y�\'��>u�l2nh�i�`ͰP���es�p��cI����Ty�U�~�o�,���ar�� �9J}�?�"L�rv:p Ctv�"Y�3_�����e�Y���7�e��0D���+GD@CGK�A9,������L?�}3j�����݇����Tޏ�)�P����>v#���H�i"|�H�.E	���!�1/$k� w��qN\[�~���SM��,_������<+��H�$�&����M�ך���P췰��2��x׬�bG�^����?�t�+eO��YN~�����fE�<����Ng�6g�/��B�Q�Vn�1�� ���F6��p��
\�@�se+7t��S@ᔊ���;��O�9q8�Q�N�5��C��tO6��C�bw�ZsGㄕ�L�>3\�fN��� B�S'�����%>{*��A���#^.f5�;�y�o��'�8]��L��v{>U��,g j��J�+����pV,������d���4����[C��<!v��.����}Z�Y~�.�*�@�(��9�5��*
iǐ���dH�`F:���A�uJ՞�m���MU�UGr������`ˈ��·{^�J�oO�i��A��1�nqPec�?t�=��፻[-�n��kM�������-���b�?���&����(Wgn�
M��ԎU�7U����	�o��Ə��D��u2���>��r�U�@�~�4,��б�L��ߗV���o�JwN�dXը�}��8q�/pk�f�a�L[H��B`(rf�$ZP&�Y�x���Q���]� Q]�+�s�P�����#6��ѣ\��D�5 g�pM6�S@��nV�_�`�9�x�@
�+y��j�1Z�U�w��ґ|�"xwכ�/-���m�X"�:`lܫH��я�֪�3�@����5�
��[Ѻ����ѷ�:eA &=O�֠8��ð��ꔦ�{�J)Vc���0�{�><:�ǒO���4.�hg	��� 
�F6�nՖ�V�vJ��:�q~�\�%t"#"����$�H��2���uV�׵c�.W�G��^!јΔq%�����)���P#�>>}��x�ܠ�.�ܔS�G�霊Pd�5t�����YpH+�X=H��=-s���U���+{ɺ��JS�� @[]��"ʨƌ.�no�`f��2D�|jA���#��	�ʎ�6�rK� �ۉ3�A`�_F�\�I��5(����r�=z��eO{e# �1%���UÔ��uԈ7刀�Zk���1�]�-�;�7S�x~�����눻Qa������2GX�%�p��٣�{1@����Ťs@�
Y�ۣ}~�X��g� ��+<\3FgM������dތ�����Kn�T��C�ѵ[x��_Ǳ�-,Wh$��Z	E�(���n q�9���a�[Vk�2g�.�]Y���\l��9����-�7�+�n���?d���c@�,��4Ȓ#N�ؾT����e-'b���_I��1UwS)��7-X\�gJ��Q�\�E��E1(�*����9ļ�{\�p0�Z��u�veS�-�gF<����v������� `n!uV��vl�!��ʶ�GNݭ��l���#	�o���V��PW�c��NSfGQ����!���n<���"Bouf����<"=���O@s��V�d�<ʄ5��kbh�WƱ�ϗ��5��I5��r�Vo����a���{(,P� �v[��[�d��ЌDf�=��߯�I�f �L6A���(�-³�� �yi����?��c3��0�:�{r��d$�7����u�l�7x~����]ϙD�8!ƔQ�Q�����w����.}�W��k+�Q	]��� �.�4(��Է�� >n	���'�n�#h����<��c�^��H��8b}���<���Ǒ,�Fx���b���3k��Y�J)V(���K�6�Y,#+J<�z��}׊����oO�n���P&��EF@��<JI��n�!y�#`�y���饰<{�	N��sv�"+�^Y��9��AIv�^��@4$�'��+8�vcI[��hv���|B8�At���ޢ��!�i~�+�|�x��f2D�cя����Hے-�Gb�����ܡ�!��:�x��^�3
�l��#������r�BQ���ڛ��V�Ʒ���F����Rh%�.��Ή7���#: u�~����Ю,�X��29����	R,b�ЛCf5L ,(��U�[�*�؝M>�֬��=ڪ�&�\�}!���z��Q`�I�،���n����G}�A��|�/I��~�"-%���}`���ɺSot���)/T0��TA�
����ϊ<,;V#r��A������l���fto��[���P鷢�WoyB����-`�v��8Gp����S�֚��դ��&���ܽ��g~9���d����4:R��c�Z�^TH���]��!�y�R��k	���5h��EH@*�2MZ;
4�H�VH��/�"���fk�!v �:�r�HC�K�{�^=߈U����+�������,GG�z���kW�ԣu\�k`��S��Q k��}d�\�shGK��"��Fb�'[��S��D?���c��8�;0tfx
�֭O�jf��]]����C�H�Y;I�m��8���lp��DrV��!���"rC��V�-��-�z�
t��xZh��S��hc�--;?��s(�;aL���M�L�:�d� _�Q���Y����D�xp١�7�m"tJ|��
H��,H�vM�xn�A��Q|k�$�W����1 "��g��_�ga7�h�ബ]�y���$9ϸ��?M@jټZ����y�o��]�� ���_wS��:�}L%��*�� ?���~�o~1��!�(��OC+��%�����xcM1
��f,kV�>X3��C��i�0�1��>T*{:T��+=Y.�a�%��E�Yc��k,��q�����L�K�F�]5"A7+��Ϲ�`��5g1�ׄ��Q6]��%�p�g�r�ϡlǥ���SO�kc--�w1�dc��4�����rt���������5ܯ���[�du�l�w����%(ߒ�U����!(<W�e0R:���\���Օa�ΟQ�J�����p���)�84��9���9�Ķ��M���.���^
�6[�.�V����ř?�$=-��4PV�w����l���X6;g�bM�����$��a�ȫhM7�!s?�oρ�A�F%ԇCY�;��(	�{�R~�'�"C�=����`�8?��%%=�{�mv����c�bH���ډ�I�9 �y�����A�]a�������ֹ���LS�[r"E�EՁ�ޔ����6���Ic�A!=�}?R���_�ߗ�E����l<NO.���U|C	sk�gP�Ε��zy��\삞��?G"o�`��pi_ֶh3��W�88֑���v؂�����wkO_�߃9SLQ��Q�_��3�[�y��<�C�غ�n��#H'g��L����Uר�	&3q
�@J�����$�cG!x���P�zƘb1��ǹf�I 4H�4��]�`��K�"P�N��������5�""c�-��/�������ف{(��S͎J+�}��*�O*�@�-�sE�P3�P�q�� ;����A�q|I���wĦ4v[¯��p�ݠ?�s\5CDph�AgA!Nc`��	����	��N�:���͎E����=z�0`�}�qW�i�3�->��M��	��9,2@����:nJ8�)��TI�r��h^!e�ﴎ�߱��� ��]�>-RM�g�����%����� Ǹ�І�A,~(��Z�b�