-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
N4/9F0+FgcInnV3I3GkAl2pJepej+wj0pLPSiDxQ+g7al8dMgiXKZUo/32Tz/JM2+CMASKLYbkcI
ySxXWv6FF8yFozKMCNCTk3pHp5uXzR6opQsF8IsgfXLEFJOuaYGN/peetOzFoWjruF3BePHLf+Om
y9gJubu8VjJWEID9AZSWckN2B0SqPNyAhZLTbBGKtzzHC3zgRsg0C0dKIe+sUajohyyx5bQus20d
redNQSEaBsDteeWLx+N1KbcsCn2w52+tqqD8Zw1Q8ecTdqF1BNn0YTDHRtpciZ5vSoRMdVe/QlS0
AYTM+dC8JxqOovzOYQirai/n0+G6COqRW2hO5A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
BAo22naef+yB1B4Njt5vtAjCAD/TE2290yBg7oKtmK/8Xz9npktMSbdmfblVaLX4NBp78LG9hooF
6fnM2c+RA04Qn/dvsW6pStyTJjwfzC5KgOmVhlfpE1ASUTE0veb5+YFrbABc2o69fEZBtpb6dj/y
VddxdcmEKI4jN6tkSmpRbU6VBLSbI3KshAJ1yijZJcQEC7QDfrneqR2EO4R0zZJZvk+kebA882Gv
xWs2T7dIuNbJh8GZt+10vi++ltmx7ohu5Xm5A/Pb0yVWR1nwOV6Z0bkTgCkZXkBkcrJagQ/T5IEn
PAqS0ELx67Alq/qRNDq9sonNw6OeWNO4eDkZhNbe6r+oPL7G7IVGDXBxPbWml070DXCSUSNOnLVF
1FjaJ4UeTz5HKQFpgXM9cZUcQ3sCCBWJ8LVnMSm97prbihbhiFkkM/V+i5fSovqmDECZcscN8xe1
zAH76IZWpkT4aQmcEot54Kt24kilg2b1GIs2tHD3354hg8WBJsrfiPUeIGkM8VYn05Xpc6oetqI4
ok4VVh/cZn9yZ/F9tao7e0kosTusSRrBYx697v+D4binHGYVP/IgRN/s2+MQwt7F30AyYsmrpvvf
3Ex47A56brerhP7QorcTzFDpdArxsEnPGEjrXzBqGMj9DjVg0b3acmSi2GNAWp2BrS+hpgWnwGCM
5PcnE6ssNC+7/K5uqnc+zeWNGf06ndcz2RIj+HHZoNaPsNZPqcSqKyOvpKyZIHZyfchNfOf4AFVX
5rmeI+RisDniX+JUAl3jlFCwg/WGojaO8aDk//WZ47OVle6nxiddFYoMuvVoqiHsoczn8slyitdo
g2+Y6Nw3UG3Tyh4sIVeLKMlJvY8L7p/1NrqqeoyNevld7HfuWL2XNANuKAwuY55JP2nWPRyOY0zM
N7PixzQgYahqovqxDY/50lzZypxIG3T3/mWFvvpunR2QY2BlG1vJXC7o6TUrO88GOrrV7PtNi0YR
XK/Gos4b7yg8IuIvfkNKorIgfma9wVUREO+3RqxiXFt8MCr8FJB8iI4B3b4mzEIDL6M80eFekOgm
sZCHeP6f1p8u14RGQnrSQzRQF6R8osmN6T1cbANINdpDxv3qBhj9xbiaTwPUJmKV3eMVXl4XgVMc
MsLPlkMeIzhUsqwro+sNwu9CxDMz/06xzWb1d2pL/mK7BRCO3h2D8iZRv1XuSW2Lbhq0bohnzbLf
sHPXpFZ/2ehz4JwROU7ftDGib9+6R2k8JBVFJzCUepIfLxGLXxWlBLl/fTHUR0xRgd58HvtycBDd
iW/XsiiJZ3hwgMKqV2PUQoEsZIRakCiY0RsOnYv/FSSgwyH0paxFUT1yb2FV/Mqe6ljb4AK47EKP
/UbXEN/2BgCEPyNK0slhWZHnaoIXjk8uNWHIXJkgZFI856qhveVa7Ij9ibCZZO/o3eWTH3giFw7e
zXiInEzkI3XpN7u4aEwlBu0sR8cFLUwKzbwZtFvlb3VVFyncdzIDnKKrAPOm4T8xWyr5EaukIL8v
SFP0Poj9LEkIa3+f1nCr6wOjhDtiWYW4WSZ/Hf/vx01SMOLB+kHhnG9yHeKdupOvVrLH9/Yrt2jI
Si7PMG2v6/EquX6+leHRgIhOO0MDR0dwLgPpGb4qFSHKjRpcw20FXFtL8vTxwSoZQ35eohWoGF84
g8D/aI66Rg4zhS3i5A3PwEk0kFjg8VG6SLoYLFofEgcw672iZDG8nBz3WizrcG/8yVuk3v27+4fr
CxbyqXkl5B99GXx7coHsvrWwQcTMl1DG78q+LWDlmF3+rghSXooVMpJ6B2dJCsCv33jtpzzTc1T1
rpoSluYQW8mqBd/np0gwghH9gs3HKaukuSsjyzOc/+vuNkF/ydnniMMb8HZ+IZNjsCCg7ZrLnt4B
OoxzbgiwdvTyDyjrb4QBcRKby76zV/tuO+N9wcfYhWuAjYf7KiDX9/smgkhLuTQSSosgAjH9QMwm
n2CFbzjmqhbcXXNXSGbDkAGQ57C4cvQOEzW41e81pcCdVvogun/aWzm46JvmNKt9eD7t0xFkKvgZ
1OMQtu1jbu+p2LWrO2+81FTNGRFbEkpYg34ikH3fki6b90LiiaxT6aDX8bSAD5I5pTQZipPJoJdH
r0yKXghKDq2BROVQaz0QY0W48QvmnL71YNpk84ozbZ02KBX7xWY5BSXF5HUaY6Lx/qafDJp+TQTa
0sdTpRLZjDyHEmuE2+JSUdu1GjgyRLcshkkx1K7jVpQfuCC+CweZ8eaVMxC/CGNy2D/HFCOOVcSr
MiSUV07+D9FYspOirXCyoCc0goOek4OHYYiTrnSyKrWntys3fXJrEDqWHLNnLQI4PuwUV9eftdI7
shQuoi+lQWeAViFql8/juW261UQJsmwFwsPGGb4dgOgivd5/x6U2CfswNK88CV2x6ZPPZiyqDBFO
AFxE58TcQxRP1HjwqkXJE54sbkfmKxWJL+gmOrT6Bkr+EE5ma38219AvmaBkRGtxmgq6hir89RZY
Db7sdCczVyZSQvq/RbHipHdGcJ9HFNBPh4diCZia51gMert+h6jthzvcfsnqI1CZg0Zr5YXB7Uca
4dfWSK5psRsZ4Xc7R8ciw28HvTRyF/z70V7IOmaB4D5JUY2SqlVmHD58mR3ZZfMbGA4k83MNg7zg
2izZISyHCYqp4I3J9Ylp8daJry3hhJNLOjVx8mO02w9UphYGJFVlBtCXz0ZwTPLjjFzqIcKru0eo
1MLv2diC/+6d21CTaWBb/oGVIo2+GpvQz0JKM3IJgHe9X3BirsGK6DwDLnRwpJgj6XPtxAyoVdav
dr7xMTn4TJt4q6IiX1fDkmh3lYtNSA/FoJl5HSBBg/ZEURGqTzb42SZbwz62u0/uLamQ4Pd0YWP2
RBHZNTmYHflPRWovswD+g13wIBrlKrmc7hcvG2tqzbtRoyZX+L4gslpcZ94BlOANZXhHEJfMwuqj
tLG8VRO3Lgv6wYBddMudae0rHMkb2P5FSAMWz+sG8+i72jhOzHMvuQXLTjHusDFIlZohhzP3C3X+
yKAD34we9ERKP2NJfWXVCJ/0Y1PRlA5Oru+imZjWXenEIpyLdkHnyjxhMbEHQif2hmOl9/5ZWS7O
fQo4y4WdkKDoP9h2nSMCFYDntnEGYOO3L2AasVvw3QI0GoLdhQyCE41fW7o/Bs/e50s5UfwrZ8uJ
nnzZcG0XhEgJqSTdocTi7AZ6pZkV9MFHmDt833c2//H1V2VFtfSUcrG6Ep/ys4rLWpUMx+C7D48Y
P1qo8j4ZuIU573xfIZFUZhoJi95K3lcbBv6e6yG3tkZN/tmVYwVVsYpvpyeJXg0uJPnzUe5YdMGU
3IYIkE4sR+DE3KQDmSwbajOEn3S0tWSPc+JftU2v3Y5JfOAb6gPHY/0FdFzYT62lGKnWhv7gGx3e
N/KD1YdyhDRLHxT8xmpnngUnjPrEX+7GP2ST7PQ3ZBLPKMFK0E1mmjOh9ApJQESJs2dJMf12/Dd3
oMYsd17zsddSAPTTHFUiZRHEWm90lhjVr/CuZyX0vcUs9qVXtsa+s2G6xZrokzRtFPuDzHbbVwA4
rZdRJJm0LEB8EeHA2DKyijRFssRjraBfGi92NJKREpwdVHbabBm1Dg2K8Yk/g2mMd3fLIM/NdYp9
9OcBvytXglo9N8QrfU+XguhEScw2H1JyYAerBX3+9j8n6SrAVgJWz8x+QOfqhyQsIWNHCYNZSkPO
F1ERA9HtTN5WfeveDeSM09h8UQ3cQHeU+VhjuikzzRa9Mm0kuNu6Wzk2SsIhYL17wWOkhfaclh/V
Vz+waxm3Tb8WoRDEv6R9U3ofsx62JuXGj5DkL0+TAUzSdANdHbkbxwm7sYeDJawjS5C7+n1WvmVM
rfnvzntADoPsIYO7VkaOM4oD8xWNgSYNw7pnvlZl2E4OFV4qsqaqESa/XY/jJnrZvJWd5SJQTqex
Pc+DzX/8HeBlhQFdTJbHEgAyaI8fwlEqJqAIyHDiyWsA6ilSdSIBBsJV7Jz0pDJlGDWx+Wg8WYze
FdbSA/juXhB9CSii+xWYY/LR6BRwHGOUfsLZWyYpRvNLCHRIo5JZ5Ttj7UZeLI2L4Zl2GsMiy4jL
m3qLNAqjH5HsftY2o5TZKAz6Y3t06Yy5iHI9qIRQQZyFhulsN8ARcVxKw8Uay73XbMMDlxKe5EFo
TZ4I+8Eps2z5QLGSslCSmXBQabJv3bLdRgvCDGiC2Aj/OrmjywYzgiVsyj3ACd7Sr3zD9tj5T28u
l39rORgtzUfuN3W9x+Zv3aGohqZ+YD7vFL2APu+mEG4Op5p0tJIvR9HWq/r5Fmvf7CgnqcwnWm2f
WsgKX4tGJPyyHS5nOSoMn1CJur+fwMf0isS2osN4waXw+5pQZI/R5hTrJbP+eXT1bUss3E+CWW4u
2sR9gITtLEs0ZO351web0BEb/A2OrI1InoXxc7NlYQnVK7zUDxUCWUlm2HoVTuD0JXqn8hLDxlaq
78i6wbtex0tNg2ICFtUq9HQ1Mp9IW/DFPIh4nDbcZ9tN4POvEBF9lUN9PBhslpHPoedlKJj6q/1a
0636dxnyDzMqb/GI7JVM9aGClhbOmq2ENDL6mUcF3bddPS5YRM8k2FImoMFb2PisB8TEbCe380cz
6KiQORnEYS2x81zn0LGi341I6kSp2TL6IBC9qtpeDlINwAcO1p/PhVUNCsX6VkGkxxXGEWEk700+
KXR5lwkQFYPEJjUk05KwmHjzx4worRo6pbJ3WOEhOBOlJY7vJk1/lLlramvGIItxqa6ROTlq67sf
aIveco/odSbjDWtaooj7ZzBn2/VuIptHLmrDMx9iBexNCZ9tkLcN7l1X9H4jD/jZFKxBvYDVxI9l
Lz0ZBGHKO3WYEhwx8pYpe+uoo4MfqFRf8Qy6UlZuFaZ9oVekD8sM7EXOEdjn0f6JFdpptDrZJ9q4
psjVbhcd/vvRM31jngePHmBs6lAVm/Ziqpq8EUVs7IjdlK3vGHKAg6MY4IJvgAN/3rjmfCbDRgWR
QWbrEg/e5SrBN2KNYLYf3eDXu3/UGGFUeotSJfDZMc9WC3WFADILXCmbIVdkCs/41Mi7Le/nn33w
14rn2ZPKr8GEpunCS05+aRAFTRQLtb1i2d+DV8iVjTc8opvcjPMtrDIJNcbppSLLvSh3pf9nM+Xu
KgD+KmJY5TR5PVT0e+cvMhh5bt0XVImkBzdXnwRJl3R7F1QEabnWqbcDB+VstiPp9O7e6lbSZPLc
d6Z31ujP5hifC3jMihDFq4I2/7LT11V25sYjpzbhHDZHHdyEP7tUD3Mese5X7BOLaXGi21lT0w9N
J8/gYTpf4llPE5KYXtQI09VX2IUJlYv2s3k972E+vpkLfIPfWFh+zLDSZJqO2hiBVON4sefxYQeo
kj8+D4Ilwr9jUVgJbRcOduTDOiAio9Dm52RCn5uluiUG2tuJK9eeRRUrnIHcEd0VVoN8G+U7r9ZS
+BBKpLMDPBBIIPvtSNrMDVAXIoV0KKQRKwCdNNI+Hkt9NSdGAZPPliZ6S7HhcOnaEdb7FEScolHO
vr41YpJUdAkcFJJh77RXasS9k2ph0k/UcAyMEefOsjV9ssHdyuUBpsCEle4xEVIE4DUiZMgkZAgd
hEFMNxmdJpMXzNqv7jF0Rj9yP91FXzj4yub7B6Mu7P1CLV39NPzSVlXk5KaB+a2QrS2R8OHc8xfW
kywG4nrNdjiEGRRjJwCK4tpE0VKQMxxboT1+zG+C4QAqm5Y1fl5Gd8lCDeLkurjC6kddj6ILGqD1
cw7bQNoaSPiV0nEUrJvpkZnqoZdz3tmrrNIslCHRYIfhk+C1YOhKV731DeNAkykoguqjRzmLkQ8u
3Mosf6Mez7wEMSUh/SdQk6uHGxZN7+YXuy20ZAvuqJtFVhf1mhGZ3MYl2YqX9lQ2GUiCDophXqxT
xxGueJkBkSJxMOnzPP/lYty+vL92ODNp3hUphg8n2VD3B5jOrOtAof637/fLSouL4R6pAbJJoeAv
dxQVn2m7N0DQ/S7uRKjNzsS5nxaRl8clTteQqudhqI5hxS9CSJE/ftqwpN/Z6/xK8vAsAu1wOgVB
kAjr3jI4WzGTmTmrG7KXnSA1leJlR6j3ca+o6+oApcn9rVZrtMkunc8/UZT37ZnlmEVI6hq1PECX
vtc7zOJNxMheXptGQs/IXsdGTyjAQbCxeJ46gmtDWiLE7DAAx6lUnUD7r65nGH4otG8+HRDz0bci
SLagdCHfMO+p4vrTobQjwOg4XsmHKH/RPTLk9XINMVC39agnIyH09xTPYC/E0qiqGjWqqVIlxA/J
yxBkifW4PCpGoxd5ALPbHXiuN4b1/4yYTxHXoDbUptg6iPAsTb0nxfs4nFMg4P5rzuDbJjozMR8M
8Fc136E+f1t52mBVXQ6j5aY+Oy9OyHsr/kYL4ZEkIi1kj1t30bA36ew97VXwSRpogGtL1xcEiiXg
Lj/1owWcaI9idxW3SPfdbRsH9sseqVhDxkSbvP7Isp9Zspg7hSdQWSBU377Gm1mZXn/3I4/9AQ1n
OJcpIERS5eIIL+XzwDODeqPe8gt4AEbb4esYiyzpqw5r5IkNfqKNtaBoYZG0ztDkuldbizkTDVWi
W3FGWaMke3nb/bsD37R6+L+bynbz64T+XyRLcuif2Y7sbpkG07mDNQqq98JHibUcKdF3ybQGIC9M
IrJ0fWX3PLNDcM8o2tcU9ZZgIPeQI1fk/voNCG1zE+zqTbEw5pDa1fj3Jvrddtyb8mp2QzCsMy7F
qt1a/6EPTdXKIbJfoNkYdRHEWNeVVu/99aDJtNhVCFexpZKeLAeDQuyExO0H03JidFWeatghFLA+
OIJeUIZIfoREov0J2le9+x6k0c06ge5GKSswYXt/l0PdmTDq99BP6lbub1y4VBqbCnaBXOGRekE6
kJNcayYAZ3a1LPrzLNqxkluyj6HU9nNkA5j5RNEJukliC3DYb5M12qhyGR/WoJfdKrB2s+GEW5Xo
SjxIjb2I9Dm1w1RMjqN1a0MQcb2KH/bAE0vKgKw8DIrz6EoELJehlPFSTyR94cFOXYhcgyRTTwk9
qfx9Mza9MX8UggafX7M+upv/n0y/Dxo7zPpkCuM85BXCgf+8PeWnMYkLLifT0Mm5k5+Ku5+C6Sx/
4XNS0Abryq3YhIG+Hog9Jd3CpzLseTimV7R0rXSkuru+h5ZE0OCjO89QaaSiynpUrzrZhJx0Ewxr
VuKSi4+G6Zy4GUdAlIjO1Vh1I8StEh78lENP+qvIdxyeFAMoYpzmrPOdqxKcSYZenjmpCLlgmfQm
ZCLZyvLP4scbvWx7mkoZhRIiNr0epRlLxvCGUCd5aB649Vj1fpx1sRSbxrlUOEN4qz/i4IinvXcD
iNI2c3OZBlfv2CerOmytGwyOT6Zavmdcidb22vl2VOqEL6Ou287/e2QNMISl6Zhax8cPhGAHVBZb
VdZy1kRLThmNHw/yNS7sgNT9iXs0mGdUI0Uo9ZxPBCtD5Ig3bFhsVhQWaZAefz0efAfyywQuvb+O
EMyMC3Zy8b9JxLcjKPnRwe0G5KjU/HEz2/cyyLvLBVrcNGtikpowgxiIVmvaxQkLwBV3QSmyWOd8
7dTxC/bjlZ7cVnxDtSFjZ4DCOZOuxiLozLQGGKbpDOA/ei497eEy79eg4NNBH9W7vY+vbt8SgqYO
E3WigPAxrb1MbdWwD7eGyzQpb6Rqvt2xdrP/8rKeLjP+4NyjsBucOEn6cfvZ1rVQURMaW3L0VkKf
/kuiRzDPvFj10vdhqyFPY2Sdl+uzG+Jt1tdd5WOw38t7aU/p4kIRfKTCIQFwogany0qQcd4roHlH
X51JDMaCWR/52tPbvzF10QVibMx0Ax51CmMrjJppfdf9qylw96ptrsLYZWBmuXTLeFrk3N/FaBUq
tDpYAq56CrHdrV3Wdk4VGyEDhMe0s3agFsoPuASVBHD7pj06cm1DpPEqa4b1uwpxW8iBgqb12oHp
vY6w5FX9Uwe+NSXwREMgB1GvQuqBlzFm8RCTR2Wzi8KptSfhwh0hBeYk63ARBIOwZcfvKBZMghd0
1ukQmax4AnaJ8WIuAYViVTzEFl9EiX9U1iq88smHY7NFj024pXBA1BbWkPfEb7hGNeb8cKuD2Yt8
hhw+kCFWAWys3bmap8i+41+2dYM88wrNMTgEKALomDLYzcQB4//+KTZPdRytXeue15ettKVsVxKi
j4UwAkHQe0tM4ho8kwfNoCmfVApSaDu/SYuZHmjN33dFzZfZBnK9Hpl5byQAMw0kEJTsjiAMaJQ+
pH9V5WWBm2/KbWBCAURVJ2+QcJXSabiuwaOpxMPctdXmNmQuqa1883jz7qRvk2cLT+xHu5maItDU
Jk5m66WUbK3Tyx4Pabv6dZ4cOgDipbneKVYNzRawR4IH3Yez5swHbISxVx8qzFRU1kmgNSDSTs43
mdH31LVZxEfPoNJ5xli34YsuVoEwXdJqmkp+qYVQ5F+IfoohaB1X9QlgkPwqs+Vd5C5mKOv8ZXox
cJbOHgZ/I+ORruEToH5Pmwp0DzcCGfnsU1mdLoP6TU2EK0vGszg03IQiuFTVF6YY9PyZK3agEQrz
KnzYRm1gHCrwhcBiJUWYuGT3q4bNVbRij3qrYiLsmNhBtkmcwAZaMb459HYntmEL7RaoHwW1C+Me
9nONdRrGt7u7C+70fQCIJOdGYIRiT93ni/H+gSspO/rdgcIrNx0hI8Vhh9v3cns/PCh9glA9Qkk4
wn2uDI9Oqtm84ixBZT/+hAhvMQ2POH+5nIAgoRLuuyKylowp43qZvFqUlb4h4Ma8rwz/isLRtBAT
jEUmMXYvHYBqMQ4virUgAeuYTrC1iz6NZ82TBwfvxR/jITjLVaChH4L2KPLPfHtDNbbxbKy4rO4K
UjEfmi8CUKdS4kqqRIz4xW3LI6pl2vvqfTd85wdhUJirQpH+WZLBCie01q1O33N5cCD9HA2BuD40
1UdCyFpQ56PXngo+PoZvRkvdSBBK2fh0WRC8bVcTtx8//KWQnjXaFBdAsbF4HN95Yu0QTDYjy8wt
LM4jwG7/20ZvRXPPL+YbgMqdrcCac7vMbWo8qSF1goiJC+8VXy3xHZNEfOvGeOx+mw/8HRV8ZShq
rHc8NkdwOqgXyVX7Y61x5hZwlXjCycZiN9/OQIiTpc4i4+pgbQ1FFUTbv2sDHQmDspcsaHK0nDrB
kMn5FuqfteSleCvaeCvDPPqLMGqKl6rrxdzHhF9/E9LsWZw6O0h914PRHi+Yb1mBMNuMlsxCcTxq
lvD4h81Yl6nEY64TXobvztpOV2fkzpwVzbWC0VbzhJa6n6fsjdEKqOpu5sza/tjBjsPpONT+ofaK
NHYP9odmJbm9A3O4yAv19+xF44Yg2W1VrFNeWM1FNox/WIbEPn+YaZ4ZUQQdYUbayb/2mU5U+Dyq
DtO+PwqaUhaYbdRP3ROLEDNaANbKHQ/2TnPyeWLaPUrhVMbAKDugQaHTjfZjzylFJIODUxORNJBb
PkQUmUBszC0c18F8IikewsPosxec35JkVkXrCHRShUrcAwA6t87bmL5q5ZWhbKS4BEME0BIEOINg
vGLVT5J2tLgvrOJA3IoGfGQqhzteLq7I+jmz0c3dajiL/GDA3FIhIxhYdX+zlmHq14WxwIKvfd/u
4p4rdx0TK6xc1ZnTOhzwqHtSKRd2cnX/IfqOh2Wdc7NocFBlknXlAJ1hQAFIi/LL4DfmYgzyJtbf
+Kv1MCbfEhxFd+Y2z5/IcxPWCCN4n1oECo0le71pOlMW06yED/n1Xve11rAIMk/ABMUdFCb1JA92
k4cHawFHGDIB50LGe/l+XfAQeq2WQuIver3YcyESSE64djfzXIyurcT7J4A2coJDsp/b9KsTpYYE
v8NG4yUHKAIx09Bzb0LJf4gc3mYfFRplEK+woHUtUlwV6alMe0GUwuDYMjoW8R1Ny02dPrGZ1psN
tgcgb6aG6KYsHLD0BqgeVvxWH3LzqGyXzuhe2q0CkBHuoL+DZ0tIXy1rJWBpjlRRRpEL+HvqFwki
l7qn/+cv0eTGPQVB1y3FcyNd7uRlC4qcuD0SeUKQQFNMy995mxOJfbNP7V21S+zzAS5w3eaeNQPs
QscOrwa4PKPN0ZRUlDjFWY9dTf+4jJX5eV3fM8cP5VeDO79liR5PuihoLp03SQ20KuHT8ALUYYxi
reNm4+v7fTtDrFCXXP0tt5E2obq7UFrTMXWbTqUZaz74wc0+u34FnQupqg92MYjzmzN8kDhqW3A3
DiAkpL/THWJBQz0vzcWGEiQ=
`protect end_protected
