��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,G�ss>ʂ�C��S��D/��mD��J���Y(�H���U��B��Z���qw0�Kǿ�(�yvE�e���e"k�^C	��?��*�#tZ�����][�5�zA�o����	�����^L�F��A�g=��М��<_C[/�
�̉2^�����|��ȿ�i�}��=,z�%\�HA&����>=��O�t��da�Fc��0�Y -� #s9�7�Uy=���[wc���(��n-,C`����Ssg��>���ybDlS�� S���x{�q�(�fLܵ+`t��pw%�u��`�B�Z��N��
΂�5tmn0"~�����F;"1Ϫ0�8�t(	�Z�x���ա~�'i��R�q��`�,�k"�`�F���v���(N�.#��:c"*�.jw%�Ծ��܎����3���e��"���˓�^I�z���s��z�P�)B/��MW灣��y�,	��@��B����Qy�-�"�pU�9׫��p��]�UN;�u����n�_��ch�Q����*kAdksP~m�L�%��*�6:9M�ѧ�&/�I;��N&%�4���n�Jx�7��\͌+fD����:2�@`��)AE1�TS�I�dʀj��G�S�DWV��>	�vz�qSL�<�x�I���t�U���p1��ӸD˘�LU��N��JI3T'@z�%䷧�E��s�b�ђe���L�y��.hm�������=t =�3}w���Ǚ�P�z�P�J	2	X|L,w�L��?9i"N����ow�e�Ok�;]�U�����s��g�p]�"��ͤJ���y�0f��Sr7���l0�k�|�� t�;�@l46�`�Χ8�`�=y���5�n�NH�C��3Y��~���z�N_{`qI+;��zf��m��-��ċ����ZF 0�R���'a?�7{ϣՊwb����sD1�TBZpD�'})�����z��4;[K���E|PF��+�e�|i�n���n�� 	���r�Jt|������-H�9�����ҭ4��_6y�kI���W�k�btf�\��T�U��-g�߈���m����'�g��I_c�$6MNF{�ˤM�3�ܘ�H��[b�[r�a�p�z�G�Ωj9N��E��+�ilP>)�=���V>{�}��$wV�5�-�QS���q��tZ�:~c��W����Þ ��W~��z g�|~����N���k�,Yg�y�pͦt����;�(x�q�b��5 ���vH`����6=�t8�����!��#�s|ӗц,i��fz�'W ET1ee�VI/!\�븙�u�qg��-R�:�%�Ƿ#ٱ0���,������-���
iL�rx��m�1����?��~G�ޕ��ҸX^����(o�@*�T��-U��/��xU
�i��5�@���f9�6��<�xXCJ�w �r^��N�.����I9�J���R{'��H�:��{�(�j���Y}ñm��SڐI�ᄺf$d��|o�M���3L+�`��m��$G[����|n���q�)I~�4Gי.�r�Y,��0H���0�������N�dCh��Ƥ�':9�d��섆�9���-�����Hn!L�V�9޲�WI��`u�;?d<��Ez�T_�ۨ�v�1��߯�8*�9���_��3� ^�������'Erz�t�CFVSHH��^G0��V��2��l�	z2�I�s�I
?��iY���
��9����BF�䑺
h����Κ�O�������/F�����K]nW�k�9�<}�$����Hz� �n�|."��6�&������c�a	��	h�-@�b�{��g4*x�۫���L���$��bY��[I����*��2m��m��˒ڥb�*B!���!C-S]A�N��J�M�1�C�IΝYG�������u��I�'"��fe�2�����\ز�=˧����Qg�����UߧQ��S�A�CZfH{Hy����P:�<@*T��Z[]��&z����%�Ҁ���G��<�/ ƯO/�U��5(κ6�*Ǽi���>.�>p��*E��HY�I��⾣os�*�j9�u�3�����P�(U���p4;8:T��e�C�@2�`��]-�z<�^ܭ�[`+���6hDRh�2��31 q��ּM�&ˠ�������Q�� �ta�hg��z�s���hZ_&����՘�:���4 2ɞ�X�i���ֲ�OH�u䊛�X�b��|�G*!Vҥu& �BIY����ܱ�����A�Z��O��+r�`D��?�X��1}�<��������	� %�Z���6�Aҿ/�2�v�
д��B�4�<�_ٙ{��-��Er�_}�4�Z��	2 x����6O�i�v�[�IY�ʫ�����T[����w��T�sc�T�6O���������Kz�eZ<Z"ݥ��e��0�N���!-L�E7��f�IG��9�w_J�FѲ��h�F�����G����ʅAu�72�w��l�� R[�@H3d�R�7������_��a����/�@4U��i��g2Mq�3])kj��"EN6����[���.��c�/����κ��5F���i�I��A]�bl�F{%�'dS@e:/�Q���7Cߺ"����\�j�&C��+ۖNO7ï(�wH�&�;�?Df���C�HXp[}Ϥ���^B���O֘�@��Q�U}��x;���H���7)-��n��)�G7��BTl�-�6�K��+��=�t����ac6��_��P�ű��9�QR����^�V��Q�l0����1��dQ�*ɔ8,v�S~K�R8%�9-V�(��,1 9DD�2����W�襎��8�Ϙe�Z6_ilAz���:=��\+r�kL��6����M�39�J <L%x��JiЗ����$���J)�cj4�1ݾ���F����Lx�Ζ�N9{l܁A�1�^M�IZgTKiX�A�*������X���5����a֋�#������E�w.7�޴�$�����LZ�j���_����9�e/&�v�òo�Q����4��?Ǌ�?c,Qp�o��D��y��!,�d9����)g�y��B���}.�XYB�"�#����������¾ɒ��\���6��;��u¨ U`\���_~��h�����)�W�ut5��4o�����*���2?\��c������'-=�ٿ�W�s��lW�};��~͙���u��hn김����r�\��|�k]	e�8�Ѽ�u{O�ّS琈_��X{b�`{��~=��GK�7�ﺾ
d��,.���[]��Q�!���]9��ߺX
=��zn"c��]{��}��:��ϫ[�����>
o��`�󒣚0H|���!�[у5m*u�X0�Y��h#T6�a?�}Q�[����O�I��O�����y�%ې!yfg��|G���JS�p<��0�X �~׬���'Gs��2�)\��3��g��ѯ����@�p`��*�[�r����R�{)=���?�s4s z2qG�d�p�H�nn4���ǖc��)�qĮN�^4($�$X�'��?�ۑ���Qr�M��V췎Þ։5����>n��e*Yk��+�Pf��TL�%WCoz��<
3?=3�2�5��/��r�mo	0���x���U�M*��j�OD<�@��<`#�g7|dH�sVx­��'�Y5��P�0	��V~Wvw��l>�C���8"���O�~��B�^�@��1~���)�=IU^�Iq�M�xl�z�h�
#_�٭_o@8�����~Ϩ4X+0Q!�-��ai���q]n�`-匵�f�W�s��x��E��6�}�y�(�7Dr�?e�G7�L�&":��k���po�p�"���5"��2O� ;���,E6,&��L�{4��fA����gn\Bh'�;��B�v��)$��l~y_��1�/]g�':�̷v��������ߟh�1C�DWi��7PX����\���M����!�U�c���ܦ4�����4�;+�5m�w"7���۩�M�9��5�|(�'5�F�p|��&�Y�Z�xg�)��-��\n�z`���@$���vVUm(oK��9���`}fH-{J~�|�������(�x�k��x�2��
�����cc+<b����t�ɕ*)d]�|}�d
�n� ɦ���׌	�je�M��iO��ɭ%��*��������3�p�(�&a�@��Q	�ޒ{�m^�-��9AWrYP, /-�a92?9^��iNSq5E�锑�,������˼��� �|#��#�%#dX� ��cE.���_���SW�Z��6���	�S�fN`h"K&�fu�5��<�*�y���k�r�s�>꾇�,5U5�iE�=ʥ�Pe�k)�����]$y`��nZ���Uz`F��G�e�h��O�̬|c����|T�VK�E�B�����LtYj�̍�t�aѯ�)���7ǗC���RN��@�q�CmA�=�|`m��n���+��`���(;�z�1�J��4�Ԇ�1b;G ��)�6��A_�J������ E���?��#�e�鴝�C��-'~�||@싴�x+Kd�vrZ�nD���,hd-��5�̤I\}�,�F��-��jz��*�H��Q�~¸<T%r)�6��#f�l�Ԡw}�=T1�x<kB���.d�^�i;,}���/r4�Qə���Ϊ���s���A����hەcB�j��`���ʧX����d�=TZv�[O�m|����65;���N|���<���<A6�r��B�%��k��8�j�����*�i�g�nH�������!b�nĄ�����맒��A�C��p(I�J{��Y����f����j�tXY��|�=�T<MQ��ak[���BY�̗`�u��C�����j��k������q"\k�`_��ME�j�fcWIޢ��Ӊ~����yZ�ME���ܰ���9�|�ٽ���qO�`�";c�%�:1B�<~"�!J0�%j�6U~�	"����n�ҏ��O��k������<]�'(a;�v9�& ږ��\&0[��/��g�_]���8?�.1��|�S��7t�0{�ж�䢊�8���nt���1�!vl�6,���9ǖh]��o�β^ �3�����L��|��Y��FM3���9�9�E"�@���O�;�b���S.p�] �{q�����E��ߺG��H��j���޼�3a��9P;�O.��2�=���3���k,�g(@���$W<Y� A��S��;�JiQ}W���(O�0�3w�'��Q7t�i�!�un�m&*8�3�B,j�Ǵ&�*h&g�p������xX�=��̑#^��d������[���$IvϚqm��QV��?o�M3V��'8|/�&-�<��7=��A�ǵ��u�&2�o�Q#
�jWG�yA���2%h�JT�1���yr��?G�A1kU�ųF���'���s�;G�����^1\5��!�"��;x��Z�nT�o8Т�n��qq���*g�0���l	�Bq$�YW�����F �&�%7��@NޜW��]蘹\�w����Wy����N	A��`��˸<�%iH�ly�s����>����>��9����z�7�'"a�>��g�V-`
��S����U��4�<@�p�⒌Fg��3�|@m>@ C�Q��y���kP�ٵ�Ǖ2��K���{�������ҷ� s��.ۅ���2�r=W0�����qp�k�K(i,i>{~�SB2�
��(VDu<Ӕ�tOݨ�5���E�4�~��+��0/F�X�D3�~�`�/��t���F3s�h;�=EnX��j`D�����F�k�w��:�JC�~�z�����rF�$^^�5|�����=�dd"z�ƭ���*��O�U(��:��p��k>����� �_�j� � JÐ�7�Z�t�ZHE��K��S��0qUI�Ϻe>�ѳ����k9, �__o_���}�f�h+戮�Ʈ��^��hY�,���%����
����y)<���Q���Hm�����M:��DO�B:q��FkmAҥ[�@L����4���BV��I�9A9������=!�N\��D�;I��:��,(�RkQ�?����>�A\]��-��hnh�$\�$��츗�oh2CrA���f2'��S��'�Ʒ�F*�p���/��p��h��b��M9�������qe�L�"�?�֞X	>MŪ}ܦ��r��#k���0�Y� ����:Q��
���$���An�L�s��`���a�'��Ih	��R���m��㹦���Q�X��ms>l�Z�S����~T�9�#��8Mܺ�W�ɸ,�����>��nB1��|ּ��#]�KL�sUM%=�l�"��P�_k��wı���z�#��~�2�sف��w�D�S�%;K�*�{�&�9����G��W �> �1�8����a�n.,	7�v�2�M��ᗜy�U쫭Av�n���ɥy�l��n����<�Ԝ�+��L\R�1(����H(�[�N���#A��_�,$�״6�7"+_��^ �����[�A��2�<XyẦ��QL�t�"D�p1�	�D�����,�ްނ�(y�x�O����?C|�l��ã�^3��V��Ub��x�T�K���q��Řp��7w�Z�I�+H�QC8b���:��~3�^�p�����JP8�M�������»n����Uc�E2S�[��)�2-�m��`��
�P����Y��p��)���)/`^F�s��i�D8���0�� �a��źǍ���E�7���v���*a�k�,��5�M�<v��P�1�hfRp��Qe���h���W^�IY�\��5��v��ȇhX{�[v���CA`�*%��CA<�mo����p����m%8ݸ�UE:Z��=����,����â��ˍ9�|(���Z5eֺ��c?%��8�A�|%��}�cc�T��o��lJ}4OB+�{,�{�vz���rJ����|��P�TE����� l��&��vF��C��c��������<'֌�D��$���E�G�(m�+�!����)u��u���bt��~; �;)z(�<��/O��3Ɗ� #eK#��
�Hi��*�ai�l�t��~���m�*�.X[�^nzLhH���	�o䠇4��^s@�������=��\;�Ǯ/eC��VA�v�Ŗ8��]k?�L��CF.��=����8��O� 	!Up�tMK-�^	��S�j�xgb�yS�- �fNqƧը"��c�~+��yAJҼR�g2l<��s�_}o-!w�VTY���)��{� �`:�������\�1�}R�̫b����z�Yk")C�@� M�	Up*�7_��F^�]J�~�`6�y�OBK=�x<�˃� "�.�h�PY�%�������
�+�:=��~