��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,`�e�(ȥ�����.���$P����)݅���Y#���X1��y���^)���Vm�e_��/H��*�ר:�n��`�V���h�U��%�H��9mL<��]�:~�'�^g�Dk7`~~�H
�93f�\�+t��z������y{ݧ�^��4�����}G�J��d�Ǝ���*����AH�N�U��̢)Vv�mh�Т$��o�X＞���}��18���C�7d(ثh����؂&L��ϫ���i�~�!��De�vV�@S��5���a��"7U� \A�I=Ί��3�ZB(5K(�}m�B�p-ڀ���}��gq	�V�����"�oA��24�(6Ys�9�?��pd07 6��K��my'����+K�7H@e  �"�W���K�J�A�î��"Z:��P-�T�V�PV��(�w�x�3��q�8�8������ʘ �v��/�(_o2�-�b-qj���X���&��S!%c�э���)+V��:�ւ��O[�{��y^z���I\&ܮi>�#j�Γ���8CK� 
�l��#��>C��D~s��U�B��7����1�R��B�hH�T�ҍ���]VM(c�7��L5z��T�v�.���������m\�`��h��Z��{ӕ.i���U����)��݈��9��o��3e�{����X$�2�CO��3��Rd1B�vf���A[�zQѯ72�Q��h���'ru{1h�bv�y	"��OFo8 ֩�`�$��K/���+��s�;���7���f#F a� A��#��<3���*���硊�e��}(��50V�2o|��s�+��T<!%��b\�>ۛ�Zt�%�q��f�ހW��LlnW�ك��ֱ�AH��TcGc7�9�;��͇�	[粶�_�$9���M
Z2i��P��'��hU�$���9���-��A��5WwE���Fk���"��@��4�H�Ģƙ[�"�*�.ߩ�vZ%�rL)�{5�����(�{7n�(Y����7��۟��<�����~��/���h�:i�Jd0���&��(A���8�K���K�#��lAk��=�i�)�0��K�p�$��'�i$L.G�%ބ�#��$� �������1��D�\D��&q�P����6�0�o��"U��n���tI��_��c�%�Fr�J�V��s�Q[!�T�{Ԅ���'�#�3M�B��_��@�͈�������*Y�G\��3E?�X�M��F#���)So/�s���ޠ�� �Vg�^*?ϕ�m��+P[#2Ұ�[�����ҿ�(4�}!����©7��y�c����P�C�X<���x�b����Sj=v��wdzљ�� ��ԙ��ø&�aN	��[�����L}�|ꜯ��!���,Ԉ�O+']�1���c 	��=�a�NW�h�At~�]��E�RYׁ�Y/�S�.��KS�gk)�y����- 8 Z4�<c�Z�L����,wr��BH��#<�j�Uf�1d@��û'	o�|Gd0�.ٱ�u�wm5e��]%u��	�(�Ҏ;�Dy/�:�G#.���M����!0�t�
�H-�i�y��GGZ�����<9�!)�10����{V����S��������])�����1�K+ ��"��0���h�ٙq�~AàR�H�QO�<��A�_G��}�X�����d�\t���7�d]@v	��+��/����6+-�y=3�pF[���kx���xA�E8wi�Ш�b(��B^�����_A��3�T��*��/qhd ���D`����ֺmUX��ʛڕ"k@�a��c۶���'����c7Ubo�ic��⛣������ݓ,=���"�Ev.�^�v땾@5���NZ;�`<�?�������`�"ܡhA����	=��0W�^��X��ٵ�&xz�)�:�����Ĵf[?�B�5�z�\�J��ځI'e��y�e헤��L])�+�s&%d�H�8��j�ю��1Bw~v�r��"��Q���7I�ey�O�2���F:�� ,`A���a%8�>7n�&"�}>幸��Ҥ�u/��:��w^1�1N���i��Q�� ���F1��l��2���0��<�8��~0~�ַd�Wkj|���$����e�k��~�r"�����s��9w��^nta���31�n�鵔&���˾n�Sx���'����lR��U�X7Po1=C�y����M�a.���b%QNڄ�$b���D�.O.�[�[��S��pX��f�����(���s�T���qBe������B��̾�+f��i��`�+gr&~�s��5&�+���;X=%�vBަ`y������Ww�!)�g����.\�E�:����9���]D���L�'h���8�G�g���}.�_�H�S ;Jҋs�o��f����W�o?c���t�'��=e/����{��}�\��c���X��7\� X)|�d���ꝭ��2=�Q��Ծ�M�	"I���3�r �����7^m�הW1wI��`�SF{!�vLe��K~���B5�5��RwL���U��+V�������ؾ���+�.���ugp�F׭��D5�U�J/��gy�
nO����xo�Kth�E2ڎ�^�@��P���!?�X�|���ڸ{��I��$(#wʀ{�4���OTUP�9�}�'�&�	�Goz�Z*�1�����6�Yi�@b��N�G�\�,A}��sjЄ��n�1��[L ��7��x��
���}�vUz{���	$6���ǭ;��v�{���}{N�+j�Z��0o��o�r��[�H��l�̶Q�K�HőH#BfP�.����K�]6��!�o�w��.�R�c���RN��n������<10�s���N�X���B���4� \,�ī���,S���k��<
�Lw�2֟շb���b߻��Z��pb�%}w��u\�D&���������kG1����!mb��!^�n�� 1FD�
c�g���T�юK��@sEJ�6J�ǯyF�v � .������Ī����e2�&�l�H��N3�$�#��mB�d��6g7ؤ.9����ҰR�HrۣX�x�=�?Y��d!��^�	2�VĤ���]
�u�A�;��26ږ���4"��dX�BR\���uo{�g
 T|I_�l�vD��P�H�>m'#ȏ��1��F�Y�鿳V������\c�����)�BV=t�PNi�"Q���L��o�0��Xw�'P�	ꍜ�to8��6�r[���]e�m��/w�D� �-O�p���g��������z��%c���q�d)�'�cp��p�^��ӄ����W:��L��@?�r�4��hܲ-��@�i{"������lt�t�mW����V��TI��/��m�J8�Yt��6!��0�	 �C�;COc\���80	�W?]�z��h�*S��v��b���w� 	�+�)�C+�b��S9�N����X���oZ3i�B�Ҏ�;�pvvu�ڊ�]b�j��5ap��4_\N�V�R�ɗ!ɀ_dؚ�"0b��Z�T8�a�>���u����ީ@�����"H�<�\X{|�d� ��G�.j�0�$�u$�:m�z3/g���W���x$p\������_~A�f�9���^`=���F�&06�4=u��t��2��B6UU��㓫뱋�����b�2���魰�wc.; l� �/�!\#�
�G�� �Y�*gQ�����7T5Rr}�����k��}RH1n�_-(��n�i�6�%D���,�ݧ�c��d��fΪm�����c.�q_���W��q˒JG�>�p��,�=��&qC`�hp���B�fG�.��(l߳6$-*�����9��x=J��2�ܴ5�x���e�Z��Ś�36���wTQ}Oy������\�Sd����Ꜵ�(߹�J���]�-����&S��K�d���m���@�)Qs���V�p(A�ݾ���z�J����ON�ܞs9�|��%�5CW�؁�e�j�*��Fi[T%�Z6e}Uyn�Qƙ#|�)A[XU�s\�H�?����¢Ja�=�
�܊���C]�g�eIg�umߙ}��wv34�"?����X�ظL���+��֬����.Bm`-i\�ˊ}�As�|���p�/O�O��L��{W�w3�����H���ʁB%��an�G�Ǣ��61k6�&����)