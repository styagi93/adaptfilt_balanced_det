// sram_access.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module sram_access (
		input  wire [20:0] bridge_input_conduit_address,     // bridge_input_conduit.address
		input  wire [1:0]  bridge_input_conduit_byte_enable, //                     .byte_enable
		input  wire        bridge_input_conduit_read,        //                     .read
		input  wire        bridge_input_conduit_write,       //                     .write
		input  wire [15:0] bridge_input_conduit_write_data,  //                     .write_data
		output wire        bridge_input_conduit_acknowledge, //                     .acknowledge
		output wire [15:0] bridge_input_conduit_read_data,   //                     .read_data
		input  wire        clk_clk,                          //                  clk.clk
		inout  wire [15:0] sram_conduit_DQ,                  //         sram_conduit.DQ
		output wire [19:0] sram_conduit_ADDR,                //                     .ADDR
		output wire        sram_conduit_LB_N,                //                     .LB_N
		output wire        sram_conduit_UB_N,                //                     .UB_N
		output wire        sram_conduit_CE_N,                //                     .CE_N
		output wire        sram_conduit_OE_N,                //                     .OE_N
		output wire        sram_conduit_WE_N                 //                     .WE_N
	);

	wire         jtag_master_master_reset_reset;                         // jtag_master:master_reset_reset -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_001:reset_in1]
	wire  [15:0] bridge_avalon_master_readdata;                          // mm_interconnect_0:bridge_avalon_master_readdata -> bridge:avalon_readdata
	wire         bridge_avalon_master_waitrequest;                       // mm_interconnect_0:bridge_avalon_master_waitrequest -> bridge:avalon_waitrequest
	wire   [1:0] bridge_avalon_master_byteenable;                        // bridge:avalon_byteenable -> mm_interconnect_0:bridge_avalon_master_byteenable
	wire         bridge_avalon_master_read;                              // bridge:avalon_read -> mm_interconnect_0:bridge_avalon_master_read
	wire  [20:0] bridge_avalon_master_address;                           // bridge:avalon_address -> mm_interconnect_0:bridge_avalon_master_address
	wire         bridge_avalon_master_write;                             // bridge:avalon_write -> mm_interconnect_0:bridge_avalon_master_write
	wire  [15:0] bridge_avalon_master_writedata;                         // bridge:avalon_writedata -> mm_interconnect_0:bridge_avalon_master_writedata
	wire  [31:0] jtag_master_master_readdata;                            // mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	wire         jtag_master_master_waitrequest;                         // mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	wire  [31:0] jtag_master_master_address;                             // jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	wire         jtag_master_master_read;                                // jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	wire   [3:0] jtag_master_master_byteenable;                          // jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	wire         jtag_master_master_readdatavalid;                       // mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	wire         jtag_master_master_write;                               // jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	wire  [31:0] jtag_master_master_writedata;                           // jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;      // sram:readdata -> mm_interconnect_0:sram_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;       // mm_interconnect_0:sram_avalon_sram_slave_address -> sram:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;          // mm_interconnect_0:sram_avalon_sram_slave_read -> sram:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;    // mm_interconnect_0:sram_avalon_sram_slave_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid; // sram:readdatavalid -> mm_interconnect_0:sram_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;         // mm_interconnect_0:sram_avalon_sram_slave_write -> sram:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;     // mm_interconnect_0:sram_avalon_sram_slave_writedata -> sram:writedata
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [bridge:reset, mm_interconnect_0:bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, sram:reset]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> jtag_master:clk_reset_reset

	sram_access_bridge bridge (
		.clk                (clk_clk),                          //                clk.clk
		.reset              (rst_controller_reset_out_reset),   //              reset.reset
		.avalon_readdata    (bridge_avalon_master_readdata),    //      avalon_master.readdata
		.avalon_waitrequest (bridge_avalon_master_waitrequest), //                   .waitrequest
		.avalon_byteenable  (bridge_avalon_master_byteenable),  //                   .byteenable
		.avalon_read        (bridge_avalon_master_read),        //                   .read
		.avalon_write       (bridge_avalon_master_write),       //                   .write
		.avalon_writedata   (bridge_avalon_master_writedata),   //                   .writedata
		.avalon_address     (bridge_avalon_master_address),     //                   .address
		.address            (bridge_input_conduit_address),     // external_interface.export
		.byte_enable        (bridge_input_conduit_byte_enable), //                   .export
		.read               (bridge_input_conduit_read),        //                   .export
		.write              (bridge_input_conduit_write),       //                   .export
		.write_data         (bridge_input_conduit_write_data),  //                   .export
		.acknowledge        (bridge_input_conduit_acknowledge), //                   .export
		.read_data          (bridge_input_conduit_read_data)    //                   .export
	);

	sram_access_jtag_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_master (
		.clk_clk              (clk_clk),                            //          clk.clk
		.clk_reset_reset      (rst_controller_001_reset_out_reset), //    clk_reset.reset
		.master_address       (jtag_master_master_address),         //       master.address
		.master_readdata      (jtag_master_master_readdata),        //             .readdata
		.master_read          (jtag_master_master_read),            //             .read
		.master_write         (jtag_master_master_write),           //             .write
		.master_writedata     (jtag_master_master_writedata),       //             .writedata
		.master_waitrequest   (jtag_master_master_waitrequest),     //             .waitrequest
		.master_readdatavalid (jtag_master_master_readdatavalid),   //             .readdatavalid
		.master_byteenable    (jtag_master_master_byteenable),      //             .byteenable
		.master_reset_reset   (jtag_master_master_reset_reset)      // master_reset.reset
	);

	sram_access_sram sram (
		.clk           (clk_clk),                                                //                clk.clk
		.reset         (rst_controller_reset_out_reset),                         //              reset.reset
		.SRAM_DQ       (sram_conduit_DQ),                                        // external_interface.export
		.SRAM_ADDR     (sram_conduit_ADDR),                                      //                   .export
		.SRAM_LB_N     (sram_conduit_LB_N),                                      //                   .export
		.SRAM_UB_N     (sram_conduit_UB_N),                                      //                   .export
		.SRAM_CE_N     (sram_conduit_CE_N),                                      //                   .export
		.SRAM_OE_N     (sram_conduit_OE_N),                                      //                   .export
		.SRAM_WE_N     (sram_conduit_WE_N),                                      //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	sram_access_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                     (clk_clk),                                                //                                   clock_clk.clk
		.bridge_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                         //          bridge_reset_reset_bridge_in_reset.reset
		.jtag_master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                         // jtag_master_clk_reset_reset_bridge_in_reset.reset
		.bridge_avalon_master_address                      (bridge_avalon_master_address),                           //                        bridge_avalon_master.address
		.bridge_avalon_master_waitrequest                  (bridge_avalon_master_waitrequest),                       //                                            .waitrequest
		.bridge_avalon_master_byteenable                   (bridge_avalon_master_byteenable),                        //                                            .byteenable
		.bridge_avalon_master_read                         (bridge_avalon_master_read),                              //                                            .read
		.bridge_avalon_master_readdata                     (bridge_avalon_master_readdata),                          //                                            .readdata
		.bridge_avalon_master_write                        (bridge_avalon_master_write),                             //                                            .write
		.bridge_avalon_master_writedata                    (bridge_avalon_master_writedata),                         //                                            .writedata
		.jtag_master_master_address                        (jtag_master_master_address),                             //                          jtag_master_master.address
		.jtag_master_master_waitrequest                    (jtag_master_master_waitrequest),                         //                                            .waitrequest
		.jtag_master_master_byteenable                     (jtag_master_master_byteenable),                          //                                            .byteenable
		.jtag_master_master_read                           (jtag_master_master_read),                                //                                            .read
		.jtag_master_master_readdata                       (jtag_master_master_readdata),                            //                                            .readdata
		.jtag_master_master_readdatavalid                  (jtag_master_master_readdatavalid),                       //                                            .readdatavalid
		.jtag_master_master_write                          (jtag_master_master_write),                               //                                            .write
		.jtag_master_master_writedata                      (jtag_master_master_writedata),                           //                                            .writedata
		.sram_avalon_sram_slave_address                    (mm_interconnect_0_sram_avalon_sram_slave_address),       //                      sram_avalon_sram_slave.address
		.sram_avalon_sram_slave_write                      (mm_interconnect_0_sram_avalon_sram_slave_write),         //                                            .write
		.sram_avalon_sram_slave_read                       (mm_interconnect_0_sram_avalon_sram_slave_read),          //                                            .read
		.sram_avalon_sram_slave_readdata                   (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                                            .readdata
		.sram_avalon_sram_slave_writedata                  (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                                            .writedata
		.sram_avalon_sram_slave_byteenable                 (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                                            .byteenable
		.sram_avalon_sram_slave_readdatavalid              (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                                            .readdatavalid
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (jtag_master_master_reset_reset), // reset_in0.reset
		.reset_in1      (jtag_master_master_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (jtag_master_master_reset_reset),     // reset_in0.reset
		.reset_in1      (jtag_master_master_reset_reset),     // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
