��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[/�������v�B�Id) |�y�r8��6���gO�=Ge֣�BΞ+A&J3����;�J�����ڟ�6��]��(�e�GQU�d��W�\��Za4�؈�a��ҧ�6#,�Q���)�
��R��!G�4���7Tzb�QA�HP�d P�P�B�4#�m�����e���!ݗ׻��0�Uy�	d��`R<����a��W�� �X��,!G��Fw�W��p�m)��dH�~mW�1E�֐��G��
��=�h�=/&�{0TBĠrR�\�ʽ(#�=���L5�/��@}fB*� |l�DY�6����9L�@�a��1��A�J��]��ԫu#��|��-���9��tf;Ȅ,:{j����V ����+Z$��j�"�]�֦4`��瑢��>�q����l���cb��>�bt*����^}P���T����?(�ȋ2��o���BF=|4<��P����(�p�Q�E�>RaO�5Ͻ}Ny�
�ERjԆ͜o�`�*D�e��T�q��&M�7�e�{�	S����>���D�c�r���QMbY��o��K�����^C-����un��ӎRn�4��{���1Y�؃UE���(�G���.��Q̋W�k6�����z���r ��Ȫ�� a*�{��	B���(�U����/D1Ć������Q���ٵ�*��x]���I�0��(|����x�5��wf�3�H��\s�0_�>�AQˣ!��08O.u�M�\q-G~r��x�y*3�`�XmJ�/��,c4j��!}�|���X|��?C5�;^�e彂���d[y�N�kt��w�5x��������o/V�B�:�a�R(~�M�3�Aߍi΅<�w汀9�nR�l wRl�a1�%CRM�B�D��7�^����e0��$��8���h��SBe�>��g�q��V��K��Bg`�d�+Ԫ��st�ñ�}P��`Z�������;�Ҋ�f,Cg���C ��X��6v*򊕝��*D��g�<����Ri@���2�.�	.y�R��g�a=PM��d��	hE�ˮС��m���r��DX'o�yy�B��#��G؞JnY��]�1R_�mU(pU��u{T�ۚz���NT�ϑ]մ\��vk�%��Ȗ��h20��Rfٵ�+����A76~AR��8E|kt_"'t�&}A��q��j�X��J����������b1zx?���*�i�����'eH�Q{� ZPQ����C,����n�O�##�0F�γ#4���"C:���SEv�#�V��Y!/�;Cɬ����kx�1~��Il�)
�2>?�f=�1���1� �k	�=�;�!E%B˒���D��_���p �8���vV[W%w��k�`m<qK���w�F{Æ�,ǆT]������"z� Ƥ��W��1�z�E
�	��.�.p���X��<V�"7P@��t��Ηi�ġ������+�`�H9<t��o���چ'����t5���ƾ
j���}Iь�<T.��H&9���.���R89��چA���s�j�>v��wy�]���H)=���H^�k�%�X�\�zL�Kg����>�&P�5}���W����-��	 ����d��;�2��p9�rC������8�Ъ)I��iۚ��(� �����J��r�֭��	V�ϗ.�y}wЈl:z���^��l(�c�P�^�&{�)�.eb|��'G7��jI�N9�'��U'׀���}7�DB��Bu�O��A��c�М�Jt*�Yҙ7!5��;�O��kQ�-�����&�[���:�$�/Q�$C_��T� �de�,��e�n��M�qճ��c�x1ҳ�u3�1�fq,�8�\⸟>��5�Z[/��į�:�H[\r��T�	ώ/K�]�ksA���]�����v�����)��~�:*�f�-�\���\f��h���˛��a{�"��g	,	$�6ƙ�����a G|��9Ls��+R�zjA�@P�y�J&j�
y����̓��� E��=�d�����p̔��Q~�T^,n�%���Ӭ�!nMJ�S<�4W��Z3O,��R��G���w򔀇���%�"�(�c?��y��M��O��x�����!��z�hi��aޘ�뻔��Q.��J'�2�v�%����r��g�/ƭޘm�4���%��M\�ޛ���>��N�p�+� ������%��-u�4i�c" S�^:Kb��g��\*���kC?	X���[�D�|S���ޚ�J&�b�����#���e�4m��Q�@���$S�y:�}'`��^kR���HȭBJ%�(����lމ��F��V�E��5��!�I�c�$}-�0u�S$��ѻ���y?e0Ҝd��B<l���e	��z��.$s�Z��#�GZax�YS�qL�>��L���R��a�L���ߤ�e�9h��n�̒kI��O�d�~m�4�S	�og$
��R�"m���x=tĲ$��~�ӈ�ZZoU��X=hD�
�77S xg�@�Q���܋?�����~�)���}�Z��W@����u��걡p��Rh�J����]��R�_ 9>b�$>�78���-��kn�x�\��";���{0�/���a�ĚLh���̒Y(MGP��_��Obӟ��{�nj�>�ں�ۯjʋeN��DnEK�s}�r�
zȁ��+�<vJ�Um��PQ����͘��9G�6��ǔE��)b���j�(>��i��
|p��3G�{�Q���N�x�!b�
с�O} ��ة�I�o�#4�]�C�o�7f
��IԆ�W9���Ъ;Nm{sNt��D^_�eԏ��U���޻�{��q��M��T�g��)h#���<Dıg����m��s��!p?o��^����3�f�2P �k���T;�2s��'ÆL���[�k�>��mF��k��4���x�SAgh�򻖔�ir�q5.���e��b�����;"%e��6� ]��\�7���f�%�.(3��DSڎ6���T�`$y�/�7C�L�Jg�g�%e�O�:����6�|�g�Ī.\��XSq&�/��}Q�]?A܍)O���W�)an�Ր��}p[zRS�䜴̱�H�W*t~�ʧ�-�`�t�Ա��5��Ɠد���Qލ��/ܽ�Lf*�TPz���-�:�S�pu�I��ܲza�M�4N�\���w��D�A������k�>ː5+�3�߻VC�]�j��qA��q*��?*�/��'w�A� ��a-ͽɒ`���-R�"��15T��@E�}g�C�Y���)���~ji؏������DC���pm����3
���6j`�Az	�� h菅ܥy0��93�F���_����S�TQg�
M)|���_�@@!uO�5϶�d=H�6#�L���J���T���EB.�`Aџ( ��iR��m���(�b�@Ơ����P������ ,�JC�U-������2���x&�$�F��,aE�O������r)��kko�X���^|&��і}9ex�w��[g�Q��&�N�������5$S�[��QlX�ՉY3�
���~�1�qw���G��
y{MT���p��ݓҀْR�{j�R'Z����n�L�U�3�R_�04i/�@���%l��/�|TS0�?�T�:53��?zr�2/W�(�F�ո�p��!6l���1@�[�p�R�	!���"�3=͵7?=�
֜F�[=��\��}C�Boh�̷�h�[nn4c�8���u�G��Wu>ݽ7F������������5�Zl.���#����tXoH��Kƺ%�-���.��Fr){�BT}y&]����$�m0.� y�[xu�׶�+��7ۻ��s��B��5��7"�W�����^N. �M�g���Wt���s���1�@]��� 5�)���~ܹP3zO���	�$�4��~����`":7$�v�M�PgE&��%>�XV�t���b�.] )�֝�Y���f�X*� ��/�+#�>=��XS�يn��6p�"$�Ġm�P�A\2�^��e&�H�"��3f�}ƈb�w?�����;GdG�_+Ga!MHTM����-�#b�Ae��w�@�*�}YOJs}�".3��Z�#|�+e ��gf��Sd��M�^x�:ٲ/� I�UmQr�S�Ǐv��̸�n�B�'�*��\�Ȍn(	1Y�u��a=�?"�g,��n����q��{Aa%��s���
�nT�4<�LU�Qy����D�>�/8ߜ�675��6��È�^)SpEC��u��|�ǐs�&Og4�YWOF��Vu��$)�y�'�� �I	dK1�r��9��dN����_��l�o��h���^[3�xB�Is�>�����A�F֡0��=)f�"3��e��X2�~������u�{�a�S0��w��
J�?��``�&��B' ����~��F�6���>��I1Sgi���[���/_�!�5j=�ZY*���ˆMi���z`ŧ]ArM�+�`qkNP;.g����X�9="r0�N�q�-+���Q����k}�W}�чk����E� 1� &����/LЗ�9�Z4��V�E|��|@�8�>�+DGt��ͅ�s/z��i�� Ā�=����]U�?x���UΕ������{�߻��_�{8��3��+̭��ӻ2��)F��v�ғ��Q�}�`P����Q�K�ᮭ���J�!/�C	4��{��9Mb�ȩ��ޚ�,�"[E��l'4������Ś
x�r���Q���k��>�&�rہ�ĕq�}X�e�p�ż�ܰϕº����Sy����"��qʰ���e<�Px1��rx7y}�D��8�`0�l0u�쭇������������yw��>�<�]t�f���ʐ����� ��0��-Xf�g�8z�BʳݶC'B�R*�{�p\�x�sVs��p�)Э���|�)��`<MOcd�B��4��`�`'`���
��$��`�5���g���C�Hm�|28��؀~ĭ��_��Y_ �0�����b�Ψo���*�N�m�z����~P�N���K�+P�^D���'��&v���<�Wt�����~z,��]S�)�4t�H��z��i�g�s
�ec^�%>�Qt\S�R�_��S��;���C5����`�49���  �1K�k`*G;n��w�k������J�?U"����~��t�k@�]�j�4�X�S��Q��4��Q�i#�uk��f�e�gG�]M�I@�ӯ��N��`n���gt�ZqT�.���=��,� $��x6�^
�S��ghщ����8ƨ�uWҒL��AI�������ŵf�����#$�RQ���\wџu��l����\,�B�C���b�
� 0��p^��Ȉ�ѕ|�)�._�s����p��%m�p�/5����#kyRАz���3 V�M�*K����]�����P�Km���tvޟ�=7E��x���kU��l��&\d�o��ҥ�CF)��L��x�z#����ǹ�]��Yl����ܒts�U\��wZ���#�;�z�K��̺�Բbg�"1�k4�+�gG8�����k�r�G�Rx��}}Е�&�BQ�~�A�ؾ����j��-�m���Am�,�06��*<o��J_�3�Pu�G^�a0s��b)���ڜ�.���'��2Q�
,	�K���,��=��3��s.e�)�Q�5����?�m���#��X1���?j� ��d�;��}?5�Jke�PiyM7�	ճ%�y]��T�#�3��r�%!����|Ҩi �
��+����=�a�h��3O����2�/�앒 XM�~��a>�~`z���9�	#��U�P��@�W�Y�^2�����e6p���޿�i��?�,"���%z;c;�u�P����]�;�����G��Q�2����T_�Lkj�j��`���q�m�WgM����
U�Y�0���{G�j�v����&�����������F?�v�= �Ȯayz�������{Y��7�x�8.G�Y3��'��6�:��z�ux�����->q�� X�4u��	�wً�֫�k��4QB�|?�k�D��/�J��Ku/^��;g���D�g;�P�fg̓�2"SH@�m��Tyu�+�KӚ֠�"@�gh�h�ݩ�ލ�o�D�jY�\�Z4E��LKȀa{�{���< ��\��`x��:Q���"(��)ϟ�"|�y/�u}wM�~����}$�L ����5�;�����W��Dj�t��5�q�JY��9�\<|)W���'�*�Z�2��mt~�1��F�ط�L�l�|�Hx].(��#�a�G��t=�/��I��N�v"��(�E1�,F-{���[}�>֖dR����c�Gh��f�H�Ț�k�_�P/�0��C�͙c��ۧ
���^6��n xr.�cyq�iP����d4߀V�0d�@��/�uP&�	A`Hf��_!����:Q��3���;��L�Jk�B�X>)f�h-�b�8�r���8(�}*��E~o�w�L�6"�x�Q[*�*Q����_(�������( Y������+D�O���s߬6�į���Z&zm�PO+�K�&�Ѧ����@�=i(i���]��g�?�i�r{oVW��ތدd��[�e���P���B�,ὠ�@� tSI�p�*I~W�F��w[�,�̩��.�<�¡�;Ň�1	m[}Z��LɈ`d]
�4dמ�%���.V��G����
��&��&���SUא��~h$(W�x�i�v�7�v�����CS������rS,Pf ��5�L>Cw:y�Q[1���3�)���Oy;�j�[Z��zG}�>�<�<p�,�����W����뱛��	^K��[��.&�z�WW�}�K�f�-��z2=��@���^�����㳗�l�5��'ӆ�a��������N&d����LB����;Z��۸���'�p���Z�Y�q/ov�,� �N92���A�'����.H��G�Z��ΧL��V�ս����B�N?�a�SW�d.��y86[�#W g?o��*��� ���e,Wʑ�
z	�F:,���V��c%�������;��\4�bך!������Ɛr27pc���K�p�r~5`��� �6�\�G��2���t;���$)XsHo����L
;
qM�w�P�BX\���/ב��3�O�ؿ�߉+S����%3-Ӟ@��6ۅ��Z�Y�yfa\=���%��-É�i��~.oළS�e������=08�C�	K<qo�*�����MN��g�Y#�3��z�Q�Yv�cL�)5r}\-�V�q��](6x�uɶ3�hE<��D|��(���T4���fiG�w}[?
U���=fi�r[G�)<[oHk�e^ғ���j=T��T����E^ަ��Ø����<?*O��l�	��t�)E����S6����3��&�^��jAs�XP��{��E��_�.���fo��q9Fsw�y�A�T3��,�(8_~��N�:��%�f@l���x��qf�1��}	g4O�c�D��`�"�׾;n� r��Ni��p; �7�����ƿ�e�6���}�:��,��q$ՅY$д�o�<c�������hw���`�k©�����bQm��P��(��QHd�a�XkAV�^r5���_��&m$W�GWW1�����(8�6b
9��Q�9o�g�?�jm<�Y:���Ř�j�|콽��Φ:�}7�.��eG��Pt���(���'�s9���a�qr�B�� ������,Ug�z�nެ�QUƌ��#oB�.�V�����R(����@��"���Un74==�u�e����N����)���3��k�n����R"���b�+RSQ��%�}��$�B�/����L��r�?d��r�٤[�A�uy^�KS���s[��R�o�\�Zv�a���ҩѢ�T\�����+�yF��T5[�-	��r��"���.F���2l��)�Mn�Y�����۵UU���ah�ğ�u����H��;	u>���$��'4JW��H���H_��
A� M�M"��'v�Bs�+�l3٠j3��G�iM]���,:�	<)�Aco�K�"�8s���6�|�*<��q9g4��4|Ç��d�����Z�r��$>��R�cP��ӓ9��˃P�vP��We���f� �D�X#�dhH� E�di�g3� Mh���i���"^%(�'��t�P=r��K�#ڧ�Z]_����J!ܾ(��F��D#�?�tǟ�a὾s���֨���9��t�S�O�Cly>�)�Q��| �{[,�P���-UKg`$ ���*�SkD=$����)=@��-��\dֳ�Z[�z��= �#�'@}"��g"+�	Ϣ�X"s�M�'U�%̢��?1`٧B��Z�O��C~���64dO��f.
F�n2N�c6Sظm���4A� ���"J0f2d�W�ڎp*�Z��^�3�����(ܥ!�#ȕ?X���7�.�/�PbI����	27s��a��&�Vn��S|4;`*#��P�}uk���"�]\_`�d�F`��Kd9�#��v��=��̗�ޥ����w�Wd�p�G�oM�N�`�T��V��Ȇͽ���k_�[���k$U�p��s!pe�;�䵫�k����~�r�wI�O{W8�w�P�Z���>,���IO�`���о��Ģ?PA���>;T����Fa�z6�1Z����aj�KI�Lg�ͱ|k�/� �> Q����&u��m�7�{�<;;[�b	��}�B<�O5}�������6�V�iGk�����qAìE�B�t��>�G���_ F�w{Wvda��e0�zm�Y�]L����K$��X�"4b(x���)S*0��-z��t�A8��_���P^�d�O71���*iї���I�'��L� $vI�� �����d��k5J^�Wԇ5�Ml'u��&�[��w��8rp�w"��Y��R��k܁`��T�N�U�*L��H�{5�mA��s���j8��xX��7��zt0R<����o����aO8�Iyf%j������w\����B��`�v�B�?����,�d��19�<���NaT;x������������.�6��oClU��:9r��$)��
 /^�^�v���Y�Tbao�i}+b����z���=���P�(#��"BJ�9�E�����j�
U��Rǔ���t	lh��K�I���V���I��pP��M~iTب��6O��-뤱y1�R���o�~+��)���>�|3�<��;Hg����Y��E[��w/PJڀ�D�,���� �2�2}�YL���`�U`6o�O@���������:���
�4s��]*ve��U��U?cHd�2Lo�/g���p��Q�����d�b"H}~��^È�w�h�V ��_��8���n��]C��i8@�-.�8+�����&f�)}�%rMZ6�Hb%�S�Q�5I�H�&|k��C��O��$ѣd��9��D{za��Uz��x9��$�t���Ta?��?�/-]B�l�A�9�-(��`��D�=�=�))K��xE��sp�u�a���Ũ��ݐ��v��y�p�)L�d�7M܄���$
��f%�t�����mCn@��U�Q��L=Z"�Z��<^�?N�g��"MTi`抛B� v��Ƿ#��v��*���uS��*�"�ۡȊ,��?Iw:��^K�D>'!JrAΔJ��W^�Q�
"�DJzR�P����z"BK�.��I������Ȅ͊R��[�u�>���:Қ�S@�@Zg`�/��ȳ��͔�ӻ�-M/3�L�p`oG}����v�_o�z�^�"H�Fe��9��9\�}��w�1�W�E�-xbG[?�Z#�{��m�y��+OЙ\h$<�h�E8|�Y!�cR��{�\@H'n�R�w�[�H["�ո�h�����@[�JPȢ!����u��LG���z��������q�ԁ�T؃��ܔ��$3ENmv��e�}�fH���� ��+9a�ա�@�T�F���RPz;���ЎX	�m��*��
�z�ƣ��K2��9�3�]!�u@���k�v6�ʊ�����ĥ�|�`/�,Z�?B��W]s��غ�^�3gByf�n�Ws<"C����zJ^ߟ.B��m���7nfCՐ6响�#��v�|���Q����ʣ[e����OvD$}-~R��i`:��:�@�!(>��;!-��I��|_��!`�q�mt��1�E�V(Ӡ	O����_5.�h2[xk� ��j0~].N���#�j`��(s�6�7�kPy.�W�S����f]�C\8-^+ą�H?�m�:�C.����,��OMIU#���c.����34'q�&��/����nNH��
ī{��t�@r[�;�"�È�/��tP��Z�G�6�M��X�J&:�n��Dwi׬���hk�Wl�c���u�� � �A�㤳62�1z�*�[U�,X�6�����_�I�F��Ӯ�P��r�rU���I���k�׀"6&h�n��~9��U��!S�����c���䗊����,Y���㸌�Ѯ�m$5�6޺�p��Ԙ �8�r�r�yS8`<�M�6W�)#�v�&B�+]��=0R�X��i���LhL̊��(��UW�/�S�@$i\�9�3���� �.��
 ir�39!(�3��@{���Ch�[�hSZf�!)�)(Z9,ԫ[�(��̔9}ʞ�B���¸f�C����9;�m[;�x��,
��t��wc��.�y�'B-	�*ݧl*��c��퍵���ɫ}�!0k��s��1�k՜��
��R��o"?Cnǟ�	nL{:���o�l���a�0O=���i�SD��4���N�����xդ���%�6����'F /%���H�Y���oJ�����9�{�9�����	�I
W�f��+�?�o������IU(-��2 A�t\��"[��d�����B�L8|FFw�S#k�;��*��_x o:�G�d�5[�p ���'q�4�V"Z��[�?E3͏A0q��ʉ�}��Bq�R��p�dЬ�l�ق( �B�05 ����� ��`�B��\:�Cf	/[&}���`P�3�z��t��)Dy�E;���sF���E�h'�����#ɘ�Y�q`��������+��\���9��E|���(_�, �Jf��E��8��|�*ǒx�ަ
|0z*�GN�d��W�3?_Ժ��~Xʨ���ϕ��I�����������F��� '5d�/�l�(��7�k��3�KHgG\��9<��6�YW�+ԣ�5ؙ%��l.��GQ�� q?�����aD]܊��D�&oKe�'���SU�g_0c�=��F��ggv�&��`k��ڣ,p� ��qЎ����M�}:�R�b!@-]�&V&�/�߽ᦝ��/��+�{��_&�l�i�De�Ǟ�n����Z�(BN�<יl�����q
�l�OWe��J���`ґ3
�2>��}N�ޯc�~A��!�R�?'lD>����w[]�����.��ڈY���PMj\�U1:���g���'�<���V9�a�oϩ�O�k�ò�t:�'m� s�|�r#��j��ȀvA������+EdIw������8��|����BXN>��P��<\4�(DHN�G�M�Ds^�+a]ěWNi.�ґs��(������يL"#π�+%	K4����,���@��N06v����S���(��Vl��J:h�4�6�B��� *m��:�g�d0M�SeSz�)^N�,v��IS������*�i(糕�|�S�b������H0��]�<J�GR�2��sL�Tz�f
�V#�8�%�i��aO|�:\|OH�	5䚥C��о����bT(��Yx�A�T����R����]�xC*vr�!E��y>���b�k@�-��C�c�l��xnTwV ��ܧXY�쟑/1�����C_bO����f�K9/���H_�?Q���j����k�
��K��i�:���1�}�p�$Ä@���;�g�M�qV��0�y�}�$T�r��$^P��d��/�TZ��TUV̻-|�����^fV�;�	~�*��,�� [H��Myο��mcm��1�]��'��,g���!�l9O}�xi-#��� !�i�5��Zb���5.�o5��I���j���\��'��/���Q��_&>��A�h@��Ggd���՜4H�/�I$�d!m�֘��A;]i}���?9�i:��-e��_�¹�kj���ES������T�rt�-o�uR>V�;B\u�F����Pd����~��{�[��33Dl{F��`Fc��:����+E?���B�AH0STMz��:��(_��Hƽv�~�������l '���>A��Nq_��o0���q�Ls�'5��:lq�H˄�I��о�6v ����t#�W�v�-���|8�_~��ti����Ei�G!���n��?K%q��mz~����D��子 ��"��~��$�1��Tt@�8Z���)��mM�sd�xC����*�S�_����s��a*��)滢�.S�����/�9�����+v��~&��,��1�2�FSl1��K
_�Ѐ�
<7���
&%�O"�s�7���*�)�b���S��ɰ��,�H=�"i�أP�ˮ�3��0� �ãj�s��?	��Uiv�<I)�t�ݙOC��B��"�4^����)T��I?2����Ɓ"��UD�u�C(��#Fp)�%~�o:Q�O��ѝ�s�X���&��5�拽�ҏ)F�z�B���>���tA}��VE���,�M�c���u�������AZ�� q1�P����b�]:h�� j��S�qV�pQ��g�K��+��s��{c�9��������o"�X�uR�q�6�͓p�{^d��fEo��C���Hh��B I���(r1���ԑ��r����zN�Ȼ�þwh8-�6{��t��{Iz
��䅉���˒�KG�?-�H [";@���UC���FN������|\VY�r�{Y`Z0�B`G��8����VP��֓ź����?{�Q��5�!Z�e)>Oc��c�tN��!I��y8m�a�V���7�^1/���ɥ��B�K�������8�G=�� ��q}>��΂R�� ���Ǩ��ހ����;������N������x��k����
�,�_�&�k���]V��G	`��B��ojz�WO{$l��PPL��|�㚚}ҧ�+})��|i-�J� 6��e�tF��2�'�	�� .G��_���Zح�eXb�f�;&a酆󀇉�O�jd�d/ѕ!�I��E#��=\n ; ��m�+�H��Ъn�.N3�K� �����>�2�2p&SB҉��o��Be�ܼL�j�v8J�]uuP��M��X_�S�kl{l��%��#�$�����D�*�c���B���eU�#D\"gg���']dS�Y���+px~s��S�R7-��������H��3�7B�;a�4��R�ݰ��r�,�nA�<��2z�V��H�=t��Bc���١j�<E���;���t2���=�w��ӷ�Y���/�o�f���b̆����-���a}�/���Lg��C�6��,̌�5�I'Q���;I3�>���M\!�\���b�pKN���G�ͪ����peR����%�w/�unP��i!�ζ���Q�EH1nv�~۶�8h����L6h���r��Jߖ�W�͕�V#8�IӆK@ַN�xȊt���J
��X�\*:�+l>A��c��=����Ǉ*<̨|O��%!�xp^��4���O]
��ȧ�C�K}2�$�L��d���'2�JAT��=H0|Jj}�+ӹ�����ӒFC+_��m���]�!�e���ʸm���D�7l5���i�A#����A|�҉��8�Yh1�g�)�fa��r�9�-�V�Q�֚rDȧ�D:8)�UJ��/���uY=)��I��ֳ`�:�ES%
��kP0J�$9t����$n'�r�08��`Q�Oa
�4�z']��?K*D���eD53 $t��3��V�E���)��9�؀T���3pd^#��c&�a��}���ı/�������Hi�W�7���XM�S#TҀ{ʑg���-�B9��Ӹ'��em5��~O����jЋ$���by�,�A�rBձ��Y��Ӭ9��v�Y����H���jw,$m�頩��I�*�Œ���e�_^&��c��
��b5�J
�-bx�W1� (�լߵ�"N��t%N"��>�\�����f�Db��1��/�g�{�M��� � ׅx�M�p�R���#rDf[��l�����0����s���P�@-��m��)H�."g�]T$B�T�V�Փ���m�����Ь�u�����X�{G�`�s)8,����"<�p*� c|�R;��V��9o/���dE�.)~���s2�|%VQ��M�6wZ�� ��#L(��#yIYxeLRBI�T�N��,���+��qs�㌥�#�b�@pF�7�9}��������k�9�â��3�d�d��Q�;�ܛ33�;~9�7�ѽrgF�0���^�D��_�zik�FT��w4������?:��+W�)3Q�	B�OxCY���2�[QP;�h5�bh�����t<��oI��	�$�D�\/ܼX�d��:�:(�!�/���N��]��"�!y$�ӧn��n%?$�?�=F}��)�������J���?O5�D��g)կ�іhB�+r�jI�#w31�a(ύ��慙���.��\7�����X�y��Xx"(378{*A3�mx�7���ux����D���`�?Z.G�㠄���dr`:У43���X����g)���H��;G�@��4{��	~�w!5,}ʙ�	���;~�W*�I�ʴ̨&׿F�_�qB�/�DGǽ�2���w�2�c�u��������BA>��p"QS�o�<x�����_FNV��Yt��
-��?%�vؒA q'K��"� �����8xDℒ$�����!J ����Ӆ/%wA+d�ܹ�b�-
˗�a�po�2"-vN���O�A�����/bF'��b���@Q��M)U9�މjD�M��}Y����{L���*�"���Q���l.�
;�eB:]\�������GTD1����o��x5�
䤂��gН������:V�JH�'LN��k�z,Y�U"��иǋ�h�|��?q�t���ؽ�W��ԓ+XA^�������TH����W�8��z��r�	|(9�p��-���g�P
�Dz9�M�h[�r$2�[�ţx�El	p44`\�r��آ�΢�#�����3�& �z4���/,��**���P忋v[�ĸT�,�]s�7�Dsd��+C{�Ǉ�C=@�p�~e� �j����ˣ�}����FaY�m��w�,�ò�ZIo+�f��15�F^�� {sj�ǼAr�
0��S�%u�F�����)2�s�5������ j\<,���W{����w?r���y]�:�Q