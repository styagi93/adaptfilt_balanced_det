
module p_sine (
	source,
	probe);	

	output	[0:0]	source;
	input	[11:0]	probe;
endmodule
