��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���d3�q	�����`�L���<ܽ�M��1�`��3>�S��0�F������en
0�@	!*�ĳ���P|��L�rH�?F�UoLΦ�d�̞Ѭ9��Y5!Ԑ��I�x��ˊu�WV`k�ȟ)�n���r�� ��G\u�9q��oUۤ��l�O;_P�ٲ��*YΝ��I~>�5e��;���z���q�\:�T���>Nǐ�S=��I�=�_���J�@��j�j�2&�����U^%"��y�� p��6�����=sF)�J�c�i�ȱR��Zz���4�1���	$zb���/`��o#�j`=4���X��ν�j[N�3W���G�Yc��ȒN��L�xlk���TY�T<� ��&*9��@c��rh�+�~�[[��rƾ�r~�z+)�L"���PJ�g���u5�MƮF:����R3� �e��/ ɥg;˅T��ZWk)�¾0�(ρ�;��W�E" {mբ��nZo�P3�l��J����G���Լ�g_{��B�ؓ� x�p���Z�^�Fja�����}�'�J�fP�̊:�'^��i)������� ,�@oϣ>��L���d/�!�;V�ۏ�"��wS^^CsH��d�ȡ��q������}��!(Oص�k�Z?��.�a�нD<�"_l�"��<��L�Z�N�6<7�p�*MQ3�8��9��.�Ev��Ub4���Go���	SP��)C�F~��O\/�z:��0��O�F[�24�Kߠ��+
dN�S܂����%4	�I��3������l��\G��'���x�b[�e\ɋ���^\d�X����b���i|3$3y-�݌�{4�,"�g�黑�����)�vKe#���29��ិU�6S��
�"�q0�� K[�Z��t� i��=z��a�/7�zZ�uF;1	Y�V4��?�j�0C���.,(%��~�٭�ղ� g�r�����Sh/1�Fyrƾx!����`�L�!P̻���ˍ�؋�����H�F�Fi���C���q�/�?4J���{�٦g&��R=	�A�ځ�CJ�:�v��n
s%�T�a���4�7�鰲!��ܫ�(O�w���nŀ���O.���eYH�LU�-��2����$�;Fȴ,_����4�#.6u����܍i|�ƁA�SH��z�Q5:�������."��B����
�T���ã��)�i�6M�g3u>a%���Xiں:?Ք��7/$��N+n\� �'*��.��F���,���>?��iO+�%\�7�U[\~�"�����<ކ�d+p|\��u��k)( <E��]]�����oa�-G���"Ƞ͝d!5�W��?"<�.�ۍ���6��b�4��Ls2Ps'W�
�͏���w|)eV�e�U���qp�99��3j ^3��G���@��+5���|)�k$c-ft���������p�q-m_��NM6�g�B���b�ˢ; ~�J���$o�4�:��V�;��S~����'��^a8���l��!���EW�?(�c;�Q�)l��A�:�������º���	��Q[X�J% k��������M�̄脯�����%��th��Y�D�I\��G>��\eDP�]7�0�3�s&���Pj�M���Δ�,1x`VZx{��Xd���mN�c3�Y���0j_�	2���^�F�:����j��v�Q���ؤm������D������S�҆�����];��bZf4�mxxݹ�9�*�������GWN�H����T�-��?sϲ��g�5���_���5��Zx�i%WLHso
t����[�,�8�C�|U}�����q_Uy9�2yIe�HpB�)eI2��,a�q"�\�밹��X�B���^�_on�}q
Ny�W�ݝ�\�ӣ!�W�3��%�!� -�Nk ����|s�QǛ~��o��O7d�F^�~�\2�c)j*vh��\�����ʙr��3�rU������dC� ����"	9��?5�sJs2X��t頽f~�*R�Uu]��ܾ��54��/�{q{*���Q�&p�\� ��	v���여����h��|���jV6���y��^L�|*V��,6�\:�����.�o��s)[m:f幎'�L��n�����<oX�b�zƞ���0�R�[eNA���m#<+=�*����Sp�,H�0��>��͝�fg �z%-Yk�R��x����=4x��e����EՍa�h$�X#�J
	{0�|�lw�����Z�8�m��0(Z��$�@.E��3�4Om����8)8E�K�3���2Hŭ{�	�L�v[�t�E��J�2�:��Y��6L�
*���s������/� �ϥҋ���D�͠���`���/���� n��`u	 w��޵@N����3���Բ�#�̙t�k�k�x�e=j�ku9�9������f�X���
�a�+0j�R,����n�R���0�D�	H0���Ɨ���6�n��s�	���&hՈ�v�+����;�ن1ը���������3��V~���U�J��b���[���L;��z�5p�۸�MA�n���7�j$��&ON\4��@yv�@;Y5f;�Ђ�؉~k��$�o�e��d��_KBj�IO�w�r�v�+zk}�	��C�j�1" �!��^��Ԅ���u�m�e�.]u�[T�hm��ל'm���-y����T��Z�y�/V��H��9�>��K)=������}�<L����t�n����U�`���=�	m���;@y��k��t.���!\ P1�����fC_�Ƽ�M