// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ewiX8vG5rmh/C23zWtH0pOmCcTgqYfrI0oLBtIGQ4nY8qev1QB4hUmZDsgWOXaTJ
CEZ/I4tBWrTkC+xmloZJ4/0SzJK1cuPVVtfDKe3TAZFvQxVwXAWPMmPn7QuiRK9O
3ThPA+AF3i3xCsinN8qZN/U7y/pGlry39nekEWeShSk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24528)
/c+y7CxayUTnsPJlgLAgK3bS850LfZG/cKrxO/w06H5ReZxD96vnnDgbqMXlewvt
lWGGEMcA9C2jhlvyf3I++AlVezhfhVNCmV0uPZ2A0e5qCTTatZOQNxvfhEj6rmkg
VHgk8qBxK70bHef5D/GhSHIarjlCGCwxPfjoRBTQmo0xzIWeWa7Ah0mItLkrQ6H/
Y7A9+Ot4vePuGfLif2uTw5ozwMlKMq75u8/F5vI4U2y2bjScvrTLYBrDYBHDF8iv
2WC1pGAgw4PUgfWwUXe9yYg0Dz3MC8mPmHlVh22eHPiZOCjTL/tzEkmzFt/ALbR2
1s++NpU8WNKcRTjPssEfx2pZxfzQjVgER1Vw/9G9Aq6IhhA1TPZY5kH14p2Hs790
7zK7YWUo4Qe+6czNJ4wmKeqwyBTEz0SsCvhNeljD0mQQlIE7OEr2QqUfrQpBQTl4
MpFREG+zxEx8EPcuttpHWFIUp0jd4w1k71yZpMGG6SnMZ7EDWGSX2oCrMbY5+rSs
qLmittoWi9jrcMwFqFoUqu9WSRRxR6LnQPml2XEFcXj5M+5I7CSkb/q2jA4pTjFM
Wlu9MLpD8y+s+U8Pp0DlI4glxxxqVuZSnS+l1lHiLomDrrMUKjgd41Iv8uY79keh
kqWNPsRGLRRo+XCuK+YI6qmbEJEiBV7sqRh+4GWUYr7OJmNpNe+lNdMqmSF/6gDI
+zT41MQ1fnS+jhjtrvRpVk79Q2y1pFTLR2OPfutueHM1xX6QGFLuHM6DdH6igwas
LkEZOJ+tv2xkJ3CewAo213ZlIYFTaRzLlLoHnKaiT4nZZCTP9sKyMOXM21RctysB
Fqe8MAXjToULDWTK7yqkPurAYQjcY7P4dSD2WtrHJy+BuVXbl/Nx0JE1bEWN3rnW
fhAW+CZ+g40Sii60NyXDXvwKOVMttmk2NIz+A2H/D5qi81ZnqB+wYvdMuSeb5xik
zQWAW6yUBwMCByeF62s+/dQ0xwKpNya/ucyLoOpLq6CziMgQ1Ukgl+dHs2uZ3FfX
flKUFWk9v8RjRSUa6Mz1GJ12NuK1DeE1a9w6miRvVQtAxpr2Z4gWNVMtozYOtNPR
CJzZqyuoyAs2PZgzzfVaR6KkhDiSUD0D4T7zoSwCTuW/ONYk77pWKfglnSx4i/D+
9JGJ5fa+zMVMcH4PCOsu5POnNnbfoxzskFbWNAfc+ADtJu6fIrBHhNWM01TufJAI
GPN9EJClaiT9UffNw4A/sxLPYp5d958hIarSWj1/2ngonQbMZxCcrijDL0rYm6me
74/CRaxWMLpHr38YNeTH3TxgAOnNFEjBlDELTWzvxsqDG1OMqIwFDWbJOGrVc4LD
lAoSuGCFL/OwZloZkiWiGdh7TjvN5Fz2U1QwHJrkYNfKHQOYD27pPM92RTv0maLD
WZT00U74gcej3t2QYUCtktalFvLbmVj8iaSvrA6Z8GInODCJQkxUIbPlToiaaB5f
+bLZYk1MSXg2u3/7zYwLvgu+7OHzmKL2W4ThQovGZZ6mycu1TIkvIYUBPQWwiLYZ
zN3lCtmdp1S6YdQtzy3UxYQZNjZLQNwSoJjA2RZEbByqVvnvV9xg8mswJQLG2qG6
XKM2y6zaNtMx7JjV5kyXAAhkLhjaAINHtnIZMi9475ZE/X3HwsvTN9UNwvbQJChK
g68gQ9k+JUAm18z9PpBxRqS2pGtAnLhGUJfr9/TRWPRUoMQ3KIRVAidasTEribxf
DFTZPY5OL/q2JeorypXWrDOGr8eopFdSY0M7F5Jjczu2NEpJRuVfgrXFH9/x7co2
9F18VOJ1sVCD6dneVAu+kroqMr9ETZx266ZiX5nE/MDRa+otzNwYObZZTsVtCk7E
V/M/CuIpSuLKaWNE5zkke8rKiBsCcC3JBM/WXc8mPr7/jbtSXnceFll1LsyV5IaU
Jpn4ftzXt3D2wjP/nDbe5o3evuwqgAqy5wa4pYyVAU/WvLOyM64ASWMpoo9Kitea
zRz36MWL9LuPfXd63e91liaTxuZ6svXyB11FG5bZ4WJgOjoRnlp2ylftVfnKcUoS
XSGz1gqQ71LfedRod/7jMnYHnPioMtWtS9fc5uXN7Rmi4MNsz6N+DqU2AiQqgL3Y
xq8ls1HKiBllf4q2h7ptQ9mDZ93ju6TAn7dS7gUYRQGTF1ia+/5Y312/q/p6FjYx
z71CIjlf+n8gvekE/Q9n1MXhPPDmT0EYY6Rc/SUdppuMGZt0oe02ZWjrYkM7EVKs
OrcdH3NVnjmEvlxOI4Ufx1hoJIlV+HL8DCAetYzEhxqm1mo+j6DfKKEH3hY/UADc
QgioGXXyaQn6GpdfEfGbJAxnHdJNQ//2o3hxPQCxyKPaMdMo/xDIlfC/CR1Pf8Y5
8my6ryf7tgMuIGnf49IGY6CmbkaESvze4J6dedlYx6qe1cnKsRJTk0zwpOT6xvnd
ZDZTnTxOR6j/lBcDMgU0ojRky3tcdvRXJ7wRGm7PjtUqg/keg+0TBm6ukO4o8Bnn
op3lORA80SbgHb7gsxzK1Ii3KpjTLpI8mwv0gf6QiRNSVmA6ibLP0lsuZgxobbka
amUH7bGlEduNozSDNpzWK+cmhQ+PjQkjW+oZS4xxEKpkD3k1bY90EPXZfOJKj28n
Dt8EMQue5+Jh/UCD2dS+cQZo2EoCZZjqyezjR8nlitwqLdmM+b2nVdHaFPZCfbTA
EktVmHFAOKuxQ4AxHO0QPZ5+qAm3sQHZY1Gt/3wioYEm53SjdRHH3Jml78pj4p5E
l2C6V8XfeXW8MyXRMPqw2SRUY3ZIsyYQeekVE9MbMij9cwwpDwZRAkhasiWv/MxF
wjQMigSAo1o6VQKfjasAI6bGF23HaVPIHUJrkM+So4rBpozk4UmGQ47QB0bNiKGo
lH7oIERMZDVe2g9FgnvE3atqw99DW7onZRnEtAcAzneXDkvRfNNIqVZGdqzWrG45
q9EWdFouciafk9U5Bi6Yq6zr9M1EroYJ7iF/dz8n+BlBeB0bqEiJBrp4Rt2TqXJe
rp/M2k97uvp9bm3F2neXa+YCU2T3meIAPxoA8jDaVhptIYNnOfFyPpLSiNwRtNfi
sCYBxtIy5ZcjVaYdHX79bNsD0TjUm0KqiycNexSGM60YMAO/rbfwbqFMd3lgFKQz
seJ2JEMbYPhCDJvYg1A4KCVIPBEHVFURNmUSrZ0WwNCgRUjn6lZquR6ooBeqAok4
L0MzSf0vGU32NEo0hRBcn7rsSUBl+vU+gdeSCt4G7wuGa3cBd8NFNEeR0zVY7kDU
DCTwMmOe1UFLuIkF6hvVHO43nZSjo8QzTs6YelAm/v6XBFZap89Sy8LCeO5hWLpl
i5qfJl/ImAir/R7kFyzpU4lutKYE+baygcST26Cib9Hz1jckzxP9Hx2xB3WDyu4o
dWSZiXSV8d5tWVJgEkSKivBch24jhd5vsE9YUgOEm79wGL0FyNi4p0SfJGFjQ3Nc
AqRzaj7H1MeNuPhhmLk8FSvuXXwSpIo8MNV/UrSjOrv4pqAjqV/bcntr7PfP9GvH
Dv+OkudKt2JAXraKZbudQ0e7ngo6ZhDHdgjZfhiMIXQqXU8K98QUpkcF1s3B5Lpn
t6MUl3j+iUnVI5iYf92xZoDqE+ssR2rB7vPpT3e+k5SSscc5k0qyHdIADcbPfUH5
7JojBMKZLSaXY56cWa8YYZZdvR0LfpX9xcW2HmZFw9golBYt7RW4SG+gLYIqr6sE
MWhZvoWS0zYnU+YvO9bYMmBxcJw82j3PIBrA0Vw0jEKhfgtiRxGKM2sEaE2Fz29H
MsLrCPGZPSOvYjKHz5DXob/KOY/yCn7SeqgPgX3D/pfeIRqymYUQFsgPADcP0XUW
yXvkkCkjPSkjcIXOn8NMiA3I/kjjKlbiahYGaPyT34PokjtuN0NL6UXTP1YNMAxk
vkdVTK6bMCar4jHx47sWWNc0LyRKbdPVjVTGHSQhN7tkyqCPR75qqOUPezOa3+3Q
+m73JcTTpYi0Xnm0pP4pR1TURHoayq9tjfJtXRFGr8MSJYHc4hAgJrvenq3A/ecG
YYbn1JNBablHjLwCYSxmCx4oYeR0mmtCa4vjfG7HGmJrNLjD//t8qF+Rlre7+Gla
AIBXSTQV2sNBuHPbFK9C40oa0lwP7MBIcN5yLscaDwxyJK0ai4RoFqaP1ytXeMfm
Kr9mgIlAIl9ruzwZCk81tdHf10WI4ovp90K3hQ5H63It+C+8++j9Hxf5jmDqlTWD
8rV58hx0jkOnYU6U/NbFTZL1sxHVKVf+dY7ibHlpmQ4Jgh0yhOlFlodbyKFKae8P
wFYHpsmyvX5JZiYNrGRI4vtNIG39A5baqNY5Y7tLjQ/IdVHLl+fQNikBV6RTfMhQ
qmkBLlHHmLU9lsYORZc8x1ITKdKsD9Th5JLpRivGPN0KJBjFiALPPpE1MDqo2Go6
A4ehWLocV0cDeeCRIeUHG85dlwzoMt5SwTWqj4C36BXk4Jo8WhgBpDIbsrKjRNoD
Kbt8YH/vpA3TRPaJEsRq42euXQHGQrFpw4JHT4nxwM061JSR2K9s7TaNhvgpFFLd
nZQvxTJ3uMG/+mD5XQrNUeRUbWYgx4nVDa6tu2UtWH6H9cCgEf4tfbQDvp73IIGl
KVYWomIyFaqzxPY3oruH6DmNxKu3EQ7p9q6SYkrounxw2yoSwkla67RgF627XIlp
NjoMdMICIHR4lwROfjSCrdtMZgRZSGPYhSKchn45VasIRWv8DesDgg15+bGqcZl3
2WW39qySCzpUIMOGL80iuDL28OqZ9jGNG766myGxxpuH5jUI7TcsPBFoNvi1Z5w9
xXcPYo4ZwCOnoo8c17Tq7uaL82IK4rVQnPOmKq16NeUIMuc+/COaqnNeCHwqMvQ6
i8wqHvhDeMsO8slhl01mKoJruXBg6Wmfzo1M1BtImPxhWEpXGeKKYRNGZocpzxZu
1uCiIfAZ5voZORR5Vulgc1sdKLk4j/0BvphK4LlT3cBY7+PBypcERLrnSQEDJCrE
JznqZc7O4CQY9lhzFlFYIUcdI8Yi6ku/g/nlsiJFDfHALzoyLbbdWlJwJlS/DpWZ
/ShRb124b6zjmA3kHJ7HFF2orXKiOd/lg0EWGuVb/xvmNDBVkZ0ixPMwZhTVTjA1
Raf588uDbmTTSnKJAcyi9nubpEbFJiLmqicCOOtyJpgI7o+UkilG1HVfkTPWF2wX
t25VnecJU0oIbohjRdhnDhuItvHUfvYEOE/NG2o5w7UGLregRpjMkXyYZjzIZKkd
OUZrMJHHY5yCYSQuRN66IT5PT77Smo/LE2MZyNbKl6mbGwNj47TIMfNQM4qHkhqc
HYAH5uuAFLSB9NtzCNaUdTmONlOG8Yw1p1nKtq3Fj+zu9sAInL+aWPPbXWkJihuo
yanGHrrCUJksjgTi2wtu6pDbMmkxEzzYHkktaHAMPD/fENe+4VxhoQ3D8JXZvabY
oUFfbACkO7jEQzHXRLnCrxuTMbFoCPLJGw91mJZ9nBMXnJNmvum3rQiVCVIefAGR
JtgxkdzF//8MuJYxNejDDmwo7LcuE4rk1R1nalkAlUCbfzC/EMUJa+DR6UyN7Ar1
J8git2MDrq1hEx1C12bqBj18jwXuV5Eb2gvkXeiAOSYtSxxPtAi6MwBBSi/c+8EC
KlceP9QNrNzoNrcS8GnIXi6D1rJhfAhGMZ6pGXVnAT+L1mzVlD4cjovHhwdqPqfG
XVxlHfKUrF0G3GPrr+ZMi4rP5DPPxsO4ej024M6nFLEUBDj9FmnYKfmxKkr8AxJ7
9PeMj3dtlVYEEc/uvav4zKVgRlX7tpXGz+1vaEt+rdMPsWlycdVBdMB8rJ/4ttxK
myHLSqwXFrigjZv4Ij0LE/njKhAeRSb7J8qNbzLoJWS0bwVjv1eYp1NmbZPvR2e9
ysKg50Cit2ygO2fYAob/iDIcTUkSczu517DpEMTJXXPsg9attW+00bIUZ07wBKar
C4ojvf62NnX82T7bYMDbrWwtvYLY4XUFdBfuo9dac3dO1AtBf+FSuM/kUmYKGpTc
ctUPfRXmNZL/fdj0Kd9XOohcmFYUhgdUA2tx5ywAqLvO2pTMvLp9VhOhoBFrmmYQ
X4TBLQUUgI9G+SWRZvBI/WXKOiw6Y6sg5+LJ1OY34hCiSTSV2vzr5OrBBgu09hbL
jbsAbG1fvaTwZBizUagbNJjoLPnyiP84D3szaG2RUk2DpyybLhyTSrrHajuomEck
kynEXPNYf/bhzXjhwBkf0Q6N0k0ZqYrlNBJdDSzF/9SsvcUMXZPp0TQf3h88VxpE
YtQtgdL2oXyzjODmO6efPpLytkw0a3mCY8Nm4w7dhy4RZZB5FnqChBAIYGiR6i6+
xICzfMqqNI+omr79RSS5BZhWNqcodgHurizmU+d7bn/Z2s09KqVnKi0O4KzJlo3o
NkMHLzXKOdqpXnra8Twg873skO4lityxpswy415EvA+3HxhKK3uF6DeuTy+cn2mz
LcCYDYXOE+A+Gqhshx+akvarvRJoMZGfkbKE+mhYHIMo6SGCwKT6KwzrfFf07GRV
9CV9Jubfkfj1AdtRFzaFbbQiqcYBTd8v35mvajKuhYviDvKXYIc87UiBSTheCoQA
J8ThxMgw00Ty7ferEF2HSeY1LoFIs5DpSUBeHLmPdvIIasT6je8LUQ5TipbIJ57C
pk1KUwl6f4nvlKyTlCMsUPf/djoQ61Lp21i/dI6WovOt0JFmroPL81Kpco5xIQSO
ZXrjvDqo/W+leDMomNgGwOptrOBcS8TfFmD+R1NIQyo66CjFzg19q2k+6JrV78sG
kGqqZwNytfDr0zSY5VqIzQCynLNIN9Da++DkcoMhRiu1Q8MNkdbyS6caZJgw/lv2
yUv8iB95s+Ficdix577sKDsYjywz+UW4oK4YLlNzl8BDFyPM6Uk7094mb89yKDSf
SvhymwctUyEAcpPsISoOTH6nTlQkpeSyVWTZX69IrkGtIqrQczdSRt5m/b/XTka9
iQrEKtEWpCnxdN+1MyjYLZ7eWYh0L/3yVJUnbKe6/oV+65Y6lvaa3uc4FO8rGZxa
ElolVlYYw/3bbHe6KZad6aLdHv3vGIbtddkAtfujo7wuT78eFVbiRevUZ8qwy556
6YfWQukMrsluPaegPUp2OsvLiIXIjN6g2RfEWiX30/PlBX8wdNFBFzznnx2cxBHP
xJMa0EPAXYkbCcov+GIeYaeL+ejSrJi1iKMYTP10pVO5LbCbKboifrjFhfrsFvgx
+jVEERKpvNbma6FM24XcBSo6+bjHPkiVZ1XromHmIGG11Iy37wHqQq7MT+TKImkX
0sidxu5WIpMtSIK3iCNqJADnPwrL83UUw3opB9pKurSEcI2B04NYvTPh5vJkxbs6
E+GUJijOv3kr1rBkYC6vt+WzgFlqG4ZEgP72xcVJqDubXEWngnnI+YgSXXKxL6Gi
5t9F3PKGwVGeWDVc2SPrW35K5hB0LO6ZNIRcEyVFRKSAk+mxSfs1dnpqlLIhUcl9
cS1eSu1PF1+NZag4jCJyx2BO4O/0DKiHOZ4pZKOuhd+yP0xejYqndY2nxCfgUYUV
25fmLbmUfMCunY9mmXhv4/hC0NCVUOiugcoCsvAR0e0fFbSymkCZczUzSQWKN41u
Illn0w78K4sG7Aw4tHKr2c6jfYGmgA7u0fmqbUKJ7qvWUnUI1y87tXsON1tXWTcl
GmF1ym4YvS9Slt8z6alKYHqPGLNGG34BX03WZyk8DXWGevgs1ku1ZA1aIrp7nH3K
bccq8zIX+8T86H5qg+X+vGFbAEYU0Ir4LkBba6KjGEf+CtWZNOiUt6YLOIZ/Rnfp
Nvngv6emER8ZeWI0eBpKeHph8GvuHmDBJIdPriKdy/qOfuNAc6mMV3BzhtnJ4xbr
Hcuh0ZvX8Bv9UUJSrotYUrdksPuBsFvwCVmuKHq/C6AYa6vxC2hKj9aCSD9a+3It
/63sPGiKue6lFyTPolnMUCWyU6QvHlbI2Hy3UpaesP7lQ9sYzP+dbfPDSj73PKcu
Ni7mmffheIAVW6U9yFxaL+Lhto1Yxu/BzmC3kHV0vcuweE1nJIHC5fBzl1kxebTo
2Tf1yxJbtM+8eRY+vrmtW7QSGJw3YbAI9zEAiBW6leFBdnIcG+zbX5bp/NxlZ/mh
IYvvBhIe5/nYvQ53GBdwzDYKoGVS+ZxYmzNnfl/CwheZtx4L3MhI3AQXZoPYPCbW
6A7JTOy9N6NE9eQ4TByfkW5oG47oITVHTVPeguBsIJdSVW5LGf6GC+ZvHYTRYQmw
MGb9LrzjVAfuMeXaerztiiUI608yYGZtNsMHdKOfqtCR8/gXmGhkkZCvpRdoXIqd
oGzxEyLmKUjKVRL39J/9MhFAp6bByei0mPtccUhnCeW3nHsc/YOfwoM4IzL1ufO0
moEup3aMViykuFbyRmubo7Yl8IYcBiksjF5QWJaz9SWWO/CdxzpZknT6CloD6qGJ
OZDm6GktIpkhaEsMVMNMcQ2H99TLNyM1xKp/gKVKBaKTdGx0ktaaAe/N1iPDAqmQ
mxskvYQZLHmdeCI84PYDESUrsY6e1hxtt8wqPLt7zUe2bCEmLjXyDou+2QqgZ1z2
XGUgigFGROuIz/tRqmi8SmmxbAfPXPskq4T/1/ydAq2rSXGPk0nbKhip59NOkDKx
kbr2vc30IzahFb9Hzm42stll2wpF3KQAsabxWBaivbh4S2BJgJK7fpiUge1VskZG
gfQUC0UbYv+AoxL6zpCJ38AhP+moAtofRVbeJ3m39TAagydqEBpmqS9D5uILGWQh
NbvSQK+0WLlJMj4Ty3vfZEDj1jFt8ONq4WW1JL8bep9sZQAsIERSpvrkhUfMSupK
ecm6gRmPTq1dwPRZeKJOSBao1nn+QKzptNZQI5bRFQ6LRKsUIBELhSs4gZZnbB+O
HIqIUkeBkVToEbC05bbmtpKB1v/DDLSyGAxyYL1At2MKaTq+G2fe1CtUiR9BRuml
o6f0jc2gQcSdXKOiMuMeB2K6+HBOJTCiiKaz2/ZJCKg9VhQUy2ltlylpRnXQChYh
NBmEaJMI9MkTQBfEgbrroJRIZ/yKYKga+kLoEMQOmu73RSMgD9EM1HWyTej94D7a
s5K2mek/PCMvqYGY45ZPjwi6hfZWJ26/x5mUGVRpvBw2tVzoO+KehxJmjoO0brqs
I33duNdMWtPbjf94smwPfBi1VL7zf28UN50c9ERTSwHNDc9lrhA9kwoELcDGM76p
pVM/CdzfKotfTCxqFFBETBqDOiv6RShabYabORN1nkb9w2d+zAW7D3H7CKR4YBnC
kCgvrkQkv0rQy7xAJ8J+5iunSWZBUjJFKh58qDhcp9y/t3IZm+b+YDys8G0Dug75
A7dgsmiRRFuKQ68q+K44emVrvoFU2qwUETHAZesSUq61wepc9C+cFui7J+9AVE0J
GXA+YzouvCxcrpDrHEYlUeku/hHKfpUelCsMn5/mIgaXV73WnOPMaOtOUpdlmKy6
38TIO6MrtpFiNWcpFUZHGjUQdv7wUocRhOwLxqVJYtowm6rmYrHkwk9nM/58ir3P
rsKK82OuIWrWuLI5+DoWEr+15DMDrll299fwNeVsIVilQL1gVerz+Hop0u83HH4o
8is2sXgWKNZR4yHSISLLBvJgIk52kMQO+RXXI0rIct8gKbpLYDBH7+R0uopPsddA
64OS9Bo2t8CbFxs/ZD0Q2OHoqyFW10BMYoHbsmrQHDr5LyQErksvwJe1sNMeK50k
r3k3W6c+77HjCTMgmZC/TGRf5/FPjZthetDvr0ZpJJino6iuyGHmQEEDCgvXKO1N
32SV8x6uN6OR9PCEKYU/z6KSe8ckOe4hTvHTa0QGY/2XKm8n8efz9S6EDzeO14ZL
RjUeaM2Ne1Ffi7K0N48fjDBXqZpCNpKyO8fs4IxEVDWMQMqCa9S45qQmqPo4Lajt
saEsFd9Cw6W0npJ6eKYwoGTXJy9TDeHzDaHNhwgW0X5es1dbKQKDByQZ+mhpMsjO
05f0xzOdYcdeQm9VpRLXajYIKbbND6Ux9/siajQ12Q2UwYk9Jjd7i6VFMY7JZV+r
F6FrIMEO+I9ww/Bj1ZM4XqeTqloNempXHfFGK8hvrEfWe/nrG+4RbruxORfXGTyR
AXbCD4HWrvjogF2RZMcy5vz10Lkj4wiFXEtbMQ7QM/KPtydesF8Cprw0LVbiWQmT
Sh4UEO9Fc0gv/SvD7GM/nAq37Lx26F8a5Ty8OKEoothG6zl5e1Veq/izj1MlAvJX
3dSIPX/6xnNqf8JQPVcegi8J56xV8s2aeFBdItLkyy4Za3ZRd6Zz1moxNQyNfsCm
sXOHz8wZ+5oP+H/+10L3zyLODSLvIU9nZPjy9E25cXk21daUzNVXSkkoADAgugzQ
uF8VGFLspN8USc5ENpDochJgxayN8lyrtVvJmeZrWOp4q5SLWvXI3JUpzSsIuZVE
NS+irc/JcIs27WE52+MXNWCWRknUDJCL4pdDpue74/G+eU39LcyVIqsmKP0vS2Wg
otoQUKAbJEYsg3Qkc2+cnnsFg5ghLCevdEkkXrb10iedo184O/ZWEJXdo5shuKjD
QyBe3ww2Qkcg7IXuqukXEvI4QisXIfPpt7Ja8inyytRJOyLFZD4rbuivWl7pGO5M
4Cmm03pkMpjMEFh/7/0MSQjFzV8ctIva6Un62/djAeA62i5mq1nurfsRWR4crbQs
Ms4osAPTpH9pBsusqccu/4pO7nA/rzDzjc/WXe45DZsWSdKXIUstzY21WqPfwGuA
1wC2cKBpLbnXxvqztnZ2AMMQmTZmcfRu5VcChXZcljQcQotjcZNt9Ab2BY+ULpvG
EONAzBG4ZFUu0RwcN31GvI3IB+Q/oznyHbBw+rYlxWpexNnNVPDI63GocLC7pBvi
zEaDImGL3HTE0YthBY+RGpIdAXZEY2xq8H94HZwwV/ENVi/zgT2pONX3BbOm7Woj
ofV6Fb5Sy9gQ/3jeT6UrfYCYnl+I6SMospkv+qw0/dKzL6DvFXN4JPfufbhp5JSC
e042k/jHUcez0hkSGvHBnP3lIr+JCRYMiOQF+JXLkrmHqqWhY3BhSY4DK5jo2Rl4
2U25iHPIINKdjFeL79XqVB0DePbVVTN1C17ltlqJ6TgsIT23Htb8cQU5S5ktDiQQ
rpiB7dVoiQopO0fFB82dhVpAXyOdP8LMsj5SbY5yisPjwbhFYjOFOUPcddgXWrDN
w49mVAGRu6qbzVgJIXHAydeJ6KUdnuD1PUtDEtUAS++NPrMe3RsQn60DVQys0LuL
dqtPTwRec7b3SrUvCDe52f9RHzgnq2Mv4FGX141kayAh6zh6SrlIevAnkZPmu69N
okt0kAX0+pEsiyzXJGiuWbKAfbdxtOj/NDV5LNIHAVlvrMg4XVa+QHVqIIKRsZlu
bS+dTaH/C1AlroRZr6XUaCe9OFbI5TREOAHhBVJsh3/f0RLvuTZvJzrFhJpa6YSB
P6Koy1qhjhjusZ/nc26Lmkqb60rycj5cS37VTMFKyS9xVOlPpNGlGDy07icxZ8Hs
TCF+DBjuVuq6r8nHC7jgjO2i71Emsnq7zKp6Fx1szfJaTkvFvuVGeDzsZvMWYLnx
XVaDfMQmsdRudt0tfMzQC9I2woCtFG0AMXlNPQi/MKBWKshD0NLnKS3OEkTbrmhq
lkrJgqy2MRdj/+xxCmaQeb26Ye3Yu2tiDZbrhjf0b8MSYEtjuvR/bipfvdddFSp7
xzjEKF1rBn6QNzjxkGV27htzCb3gf5JAvJK8dCREejuGKvhk1xvodv2L2UVWM4xd
v/Kpc0rbDIil90/oKM4P+UpeLxsHrON58RaK82KnZfgf70aD5F6Ik/JRyHa4zI7O
ObpZA95e4Sr1Q/Rz5TzIXg8vlhrFKWDrFARYrqXdAjP1xnpSKj4Hyb764M+eOuoX
e4IW4THZjj80K00w4Mbo4YhvKsCVUL9dN3qchElHvMMZRsQySWnz7sWxw/dyVyU7
SSb389FoUd2qQ7z+l6nMhZbiPSK6kRiDfu8vEw9ge60NBmFyvCl18RUAEPVOwYdM
Wd0QFynVrhhjZW0ouBbeKzI2K7Of69qers+cxAnjS4vlVCqtooU8SFdVmDcGDE/g
/W8E1zUS2bajXSZpj0yts3+UBKwCFfsn+bxKvVUBxgd+A3lv4A6dRuh6Sxgvu5On
sQHVkGINlG4Xcj21EN7PZfnP5kOPIqC/D9ucb2H4RmhauTHjScy2oG36jrZdgh5Y
BEZzDEAR6PBwHLVOfmwyFaoeaf1hyCnCedWOTVbQiPLu76Mbo7e3gLwpFP8NPsre
BArgj8jQq4iY4EMMDu1AH1mmHqRaOGP/ye6sMi+o48OGB9/euKU+wSR0J8DNr/9S
mSK9Ha28y2ECe/LJruGyInNFSks29+O7w/NWGpDhqy04oiMrJ578LVAcKf7yNTz0
HnAS8/q/aQkwSfAifpdlBEi2EZs1r1D//uQrSj62YlomBA4bRkqXDFXZC4Ujzh+2
yx/IT0C4ZlssMwB957LfVAEUS+W/RnKnrZqiyzk/E9HN+mg6kGTcv/Fx6oxcAaBr
Yjhn3TXdBAQCWBJFkN8IHW9U/N7Xnum4/75otc0LI3dsGbOaA4HruNzYVTjGhNDH
IUsGfVRps1GCzXk+4bFgb2fhjAEI5DRg46dlmosk8Z/f4cYDSC1Y336xvR+O98aa
tNpdOz5Df2au8/mG9jXm4FB/mlTPE5puzmLSL1ioLX4rVz7DVNhhoHbYsNdtr0eb
gZznTLwt0H6EvCHaLsEbEYRHqm8UYXF6uwMIflQjwPQWlBVihMejc7Nn6LmKjE8+
w//c8gCQ3OB+vw5HcwirLlpGHeT2LFZA/O3F9LLNkj/FllI6BOh2bIKaOUZyWpz3
HPug6vsz2m5i0i1KErddUmxzBp1JqkBMXiRFJ33DD6Hzlv13CxszBuBpqGcK9DPH
NkXSecQo0g/wE6TXEqv63xkLAyx3ODeAlampOVg3wolUp3FJBvqjVvnLnlkpBqNJ
0RqpfTjEybSbLKS1ebKWuimvBrMFoteJejmZt0RtzCVK5VLYDJXG/WeOTHhxsCHv
pBM/fKbxfz24wXutrkFbm3uG3C5NupFnJofjbcWtm3MxswWX9Zo5Yy3cj3QHAR4F
PIU88N7ot5WAOj6JqbVbG0Bkf3CELM3KdTxWzOy1tt3mMCsazRYwi1Ytp66cYN91
yTHVXJI5FPQMV2szyUnqpNA+ddNzwgUZi0oHLcra31PXkRVTONHVTO4JFxiBXZu3
3wn2z2kUg8l4BAfmZl+QlcpM62y9a6GF0LBpFoHUiqkUdsJt99+nIU/ffmsrPrV9
u95qi6BY6dP/imfnI3WJLR4nSIJBJQ4CqAM0oJ0q6w5gAGXLsPTpgulGc43qyxT4
0f4nuEv/+1nT4O7SGjnWCp07A8oL2/2BrDj6YDjfRk9VQJItewTV2jAlQYXI40g3
peQkNpEhyePyR/EK2lIcJnpfKRAKmYWMOTBncKHiXQ5R2KqOogCLIvhB5gu+4K42
73MGFdF8ku9fLwi3uy51HSHDGOq6KpKxgrIfLf8uBk6uxwy/JB+ggdRnCtPqN/Tk
KFEIzbLrkqVklOqEBmYqCbORhkJouvgmcQ4jpCBDpJr1lPmaRuzyC1Nri5dOFLbu
OaqfD8Kw6cRd1xC4/04IXrz/tSm7beLAqjYklF84ItbqHzjTpPTrYnohmwrYGIDd
Mvnwhj3o3XqNWVV1wmz1KY3JWb0IFG2x45HPtYgs0/a86jZU2K/UkOIA2h/BXvnW
wB/6uNi6jYMSgkUZgNzgbY1bU3gkgb9OJJUenJOqc9IBh+S6RV7oCS72y8FdROTg
PzPFlyZ6B2RgVfV/1Kc31TSgjaXcu7hemx/Y4t0vfMXRSHVzUiDtmQqmJXrDujVC
cDHFtPf42qauKsbBRzuqybcn7Kga295+VhATx7EezTwQhTEQSNRy3+Ms4v8ykY6U
Ho0flFI51vRHknMnlM5a+8pO8FRaxIh3FVfjnKersvQfpjeCSx9rsLvmN5/OIOIH
uh9t4oRJ4+/ojOlnVSD93lVmJSpBeZvOEd0WV5fj+16p5WTeRnPVLw1blbc74RLT
WGFNuuY/jadtr6Gap10DWyR/B7MrujnoLCPb9j/mYYGErsGERo7EotiWj+x/XHoQ
Qd0Sdv0mJBXFRUt9tdff3/KnSFhZYmopWmQmz7MhMxpx0SxS3XA/DYQb2gr0fIJp
MbWMuQqWk7P/OTj4hnXmV/6+SjRU/mb/Se0Uvi6BLsI5BhC7Nf7w3B10iFDTmQIS
oDwFdSPJUOoCr/A0Xt33C6FsXiyxdDE6q82zXURBpVf7sMqxoNlLXXTw5d2+bmjl
EdQ2zY6txEV6vor69ELbuoua+60fATrymlQ4ph47c2ngfi6eQ/otazx4S0PqG8MJ
UulpGoYoNp4b6mOSiQhCPkNXqlOSEftZl9ideuR0Wm3V/EPL2IslhbHUJujhpmoZ
d8b2bfVB/vFY697mT44yqi9jVBp/egMrAfPgQ8avCaTZozoKBZR2x7M89lPXeNYE
QsYIK7rgD59aIDM6Y+bWTV9/gQ/ucSU/uckuEJtOnLNVbL8FjBWrjvshVjmoUKSm
tuY5C5B8VcmiI/7bz6ukAUTzmRx/gJGZ0Lffuk/GMNtxGHfJusKxOxrmIdyEsDG4
WJy6jy2pCLSx4ZMYoHap6VwH1Vwjl432DuDj6L0KmCjwbRjdAZbZ1vvxB1KoVdYO
oLvAJwkWqbbNiV/LRkN+yz8psljhAJAtDZdCI27f+S32jnA7lI2YaseY49cp37p9
bU8vIEnO6ZFZubY4QyN0yeVPM1yFbGfyA8WyBNA1W0xvs8/Oti9JmbMz+rWpQS9m
twbYfSUWmtxdjpQEpvwSR1j3kUTAKUSexOmETwN0C+tpB0osb+jrnwDXC2fH7kG3
vff+B1kmqQrq1jqyAC/DMSImxVEAh1g7sgM/z/62H5I0g9yr85bDXlxg7JLKRJ+F
Qzvef8ET7IW8h2tOC+WDdcfKhvK0WDByx+8Z7FzfsmyegRGddIf5bCZ9kMnZNJNC
QDq/OBdk2sjMm3nK+f0HIqlVwt0q6iJjuG/SPJefUvVq5EKjcLTmeJjx0HOQ6Ii0
vBI3gCqPtBzrnxEJGQANB4196R4hYbgsTHmiOW7Kp2kBysOPahI873z5GOlvTxrn
XDMxA5+mUS27ffx8clwNg5zw+ZqIbvgKJD51KDrNumLj/TbBS1wKvdQx/19jXgPD
IMxA+6+jCKY2oHsu6QXKnMQrT8mP0Yn73/AI/tsWkQWyNwhd76Z5OCBRS25Pqu1c
AOO2pw8l7QNnd0rpdQ5hCtbgYxRm4kwFiuBnyEdMr3r6RiJWCbEcgGZQznqqB16F
7F/XoxtHFZKCAi9Vv6I7C4iOBqUL+aKOqlYUXSNSclcXVrkwzyNqxJQaH+slMAj/
BQO+McZiE/zs+OnHjREMvTAKamcBr+Z8WH79Vk6zLtEFPAoKaeub47lSEuIIx5rM
ryNERXpM9bbxDX5u/m11Nwlg7m8jmcHvdpCDg4i3xmzwEhzmROJXCQBuThm+UIcg
2IIGz0DQuh07Iha5Ri1JGEdUF28KtJDTuxZgGc9s2rQDlI4Ae+iyqFM2tBQ8qo6P
2xPkNk99kUAIzxJOldpA2XciaS9T9/K+4OP78SiMDFQWuNj20DWrknz8XEZh3MDV
yoLUc8AcKJMKCfCL8Ze1+vm2YDbcOkXg7U3Z4GTpBAKHtcrnCeCGC1bJ/BiKTjQ/
RoUVJTmI6pxgLgOSnVRJvkrF3nr7MFwmLX+ChN6LTBASGtAaPssAr5I7tIfbSoUC
UGoLPUOUMWgTmKcIlbCXqMifoIEkTT+pqwETG7TLS2tolMhBTNdSM3vLN+yNKtc5
9PX/B+dyR3VFuCUWHYiEY8hC9EVJS0Dp1n6PErCt6w+36nCi1HmxaYiqeIIqAMsW
U3tIsz2nTjh66a1M9NzV64aanWHpQJyGUcQVSF0/SrtE0aM/xNvwRq/sV3IQOCkS
zgSiv31Ee+2j5FqFrxPXrBZqhGkzQ6Bmfy4hP8CsBwQ4eZb8DnQPE/uuOKAvSPEp
DjB+YcV0PN/Pp0x2SeGACjJnoI5ej6uOHVbNdDqsy7MbgPyqEKdRdWpvNQd1sv66
mCnvCFo8onYk/FVMN0M7N4GCq+++uKGZz+Ef368WcZoV0sQl4HGk2PplkHAMJp+f
0vJFHhfY21fex9qsC5HxHi1j3CSJeeUTPqZY1Y5Qgeqijc+slu8UZ13G60kmqfFu
epTzGECPECDiK3zhuI5idoIzwkD9D/tx5hELcoGvhrZqzQa7tBglfy+OK0+lCMxg
rxsA6PJ4D6u5sVXPIbLMC2VJ7oVfJQTim7vWloDdB4YHwuLZx2B/rmBuigdgyn9y
Z/xLVyM6Yc5LEpEWLG8wHgQMegp70i/AqxDnUgdpHW3K4AcmqcxYUYGgOlev91d3
grdUC6iqCd2ASTWGlQQZmPJBHHDnviAwUbEIBp3LsU8qOFaLLKd3ureEDzk+GXvj
3Kv1mITz7a/UJ6JpN0eEEJTWQtnyfBGcwfrJJA3A/+igieHOS5DkhXGVQ2MPGjAH
6moGlDUhPgLTRQOK4wEltCwTMIrKojnKkzie+Q/fxtRmdn6Grb7UIHGVkva8Rk/W
siqioytvjbxQk7TsQILNzNjFSiQZ4ZyZB3TlebKF6ygl1rw4NGPI1iYITiQ9qpmq
IUCbCO6nUHlozduw5x5mkfDsBCp2ztSHYKfmDHuDeoKkRtI341j2uRu/EXIDoVbp
/s3JyLNXrqIi/q1FQh3rwr5cWbOmgbIEGl9/crtem0U7ssJLN8CHwc6VKvUHEUym
qxrasWK4GThXwjiHifjoC8CChnoLCJvZ48pGasebUGUyeQUj7ScWVXSh2rUl7VQo
Wapr8ubypI4yDfCV6JLBatAiwianl7xrDTQQGJQqpAF3rVgpD6D3XdZuuJAlddRI
vGUfDEU5LeT6IaZ6yBBI4USwjny7WaAQ+hMxkiErZYDdyVsGhnUqouLsCSVv/WYp
2hYcPc9xEwDxx4seHoqbGWDTz4BrvIMiWanil1JgllTyrWxuUomZnO6AayXF25ha
TSlXUyQ6DLOoulyROJMYGQaofBTWfxsbHEWhyY7gk84GelL37Fx25UUkOO1cOXoD
3AyuToEf5p1Szts5aVMuDfOZ4vLHI1GRFKlF8/JqKeHOINVJ2zfdPtT7KveVdpnr
2MjZUQY0Vc17h0+lG7uQlf8GbonXxDu+H6Ds7nu/Ir/BI3zpAo3zes5KHcjJ18F/
bkgSBxOmHwg/1qyhKiowdIxydLTHIJoD3objaJfAGorrZ1p8lEpbV1k6ICnEXZr0
3BmbpBVgn0jQSlQnMuBEIAd4xh4+kBeaaY+xws+NJqzbkFDX2kGv+2MAYwB+VdBa
nce/G7eJBv6j9FI6GC84u+jckJpctNOn2m+mMYHhMNyP3P7X76Nzq8J0nmyauNZ2
KHNDI/cJtK3yquNyFAqT5KkbWyLBOLkWL6JwHtYqYmhWPlTqZOGCkMjDgYPADUEw
kzWLwTKVSY5OpyQDhBppRqoHvbrZc3lNEt2Z1QVGHMy1xPMODfLZSBuyQYAFPhOU
jby7teNX7hbvCHgdZPbHX4QgS3Pq+DqHs4kkzOun7KLRl/2UXgMbOXnLyDT9rJeO
vZqem0Wqgi1I4KBPIvqecxJvVxDg+JnZJXwzCxECwtQh4oycCNmeQlWUgD+h7gwp
ZK9/jW3CB/DYNEfGYf3M7SVvI0Q8D5F/cAFPlMvcz0ZSqK2llIyo+sxUDj3MeUZz
53zfygCfXt38iyzGHMNoNfqU65Df+yrIJEinbHANSTA+VGF18YkXoMvkylZ2N21q
UHMrBeBvpYXFpHEE9L8+XXd9f6riubIodUV2yxNKuTRV3UEXwK24s0ngRRv9b12y
Uj9xxrDTIQ1po+wOtdShSotoY/v6FsZasYPkLqajoVpf97uC78LOjXlTAi7+OBqL
heOfMI+hdg1XGl4+sAYB9fjbfN+c0x9U8qjVSsuj7ah9M/EOFmhWDZ8eKLbNzL5i
6AmlxXSfzacoLSLfzPUDsJ1R4E2WiTfwSafWWYJ1LapfD7TIKye3M0j67O1j3Zj4
AmQGeCEjW5OxfKXif539oxeAK9RtokjSBmG2yGFSxudH7+ZGrkN7fnBnoK6A8H+G
aafbAW0Q9jE1CUlDeQbPJPWza4vrWvnOolIb/cOSNAlHUQ6ZLnS9zX4YVmCezUcD
gcDNH96/ZBs03PmqS6lc2oLMXyQzb6v5q3GCAGR5J8Oo/K4Y9Rt9vs6dlHXYx1Ah
a9f1i8+Jm2AA1MieGFFQMje5foD2UlbWuAruHPkRKM+g0DNp3LOTZTFAlH2dBq2J
SxUwMpLxNJdY6sNLypHZI10xsamHkbfwW09Hk1V45QsFGEgZdZyHrnzVac2Qqj/C
u8D66YE0vBWiFsbbwtH+qRH458ncNbNDM/uglv57S5nX5M4ttCOgZpUxpPwibIxE
p5WeHtt78WwCSizHHhsqrG0qdlcl/Ip9Lbt5yuIXuBfKo+/UJTZPzJUZ9zM7Hpw/
dZZHvr7sIv0jYuutES/KMJWnzYlK0lRGe8tbCoq6n84fmCdEk6hwgDYVHZLEqBuw
O9zdmxi6xAew+9xjoLYx4TNBczZL7jgNOUosDDXITWXAbQB6j7AzYno1IX/cJXg6
4LOpLyklp7e2azcEwuGDRgKBtUdeDF9LBM0UaGIeIcUcL8S7SdcN/2S2Frp7UYZP
oAglc9VtuF3IM0EuzvmxdJOrjPynjZvQK+nevh/jOTeTai0teKPLHiqUUi7vgi/o
gpeWSeAv0450F7e21N/FzlIsUL2oMWu0jEy9YGpDG57MXBzrYPRLY95VkLxgglX+
zkwKf1PR0XDIdOUbQ5T6GsxaRUXt+EBaVA7cbneahDLjzmN9cKrmlVPjkLJStrKI
wffJhgJsCpJ/WkbyubUYJOynWEkGkD0L9dJ3AsuMJdrNR9c3AbZBrwpKoqAEv5MJ
HaQBUL9EqR8GFmiSB9ardc1SnfxM8t2xHmuQB9ZXi4nqUjMJQq/B1TNbZ+r57uam
8sqF2LWG5tkjS0vleUSa0OuUQs9/PttJVr1/tjfPW419AMIccyU1v8JF79NJS/uE
j5SW3gVingfeM1d3vtpD/zjXbwvDHInUYRMufhfxa8P1X/Y72s8ZkOV22Kq2ZrfM
XIFy/QoWvm4hWiTg7QObG0a3Vn/ffwL0BrDVhPO/2PfVP7l8SJV9mxCGgV5TATba
G4DyasXhmU+In0QNiy/D9R1iQ38fLX+pfGCus+M3KyjLdRr3DWcgljFvUh7EWp21
9rALzbSdxlBWz7IFAv0xAomOQs6kjII1cf8827TlqVsURGwpBP0Qtjsr0T2XSvpg
hVY4fdICiwaN3zi5SVIaftMR5pz01T5B1I2x+HalexucN3k7LodlRAQ9GR1TcmU+
hB9+xJJZCnFhl7yBjtuj37lMYDyv1/tNLv8VbJvEzXXz22+s1DFTJUHSafeMYtAI
ARgO4hNxOHcGwOCf57RVxrznZCnd/vQfGPrf7v8EoDGMaUZJTezNZOu4iD1TyyS+
F/MxahBSSvxXVr/fTPmKJhn33lfoxmeNfG027zPZbpPgOnXfK9YFWjMpxfCZ8PKK
RMnhPvNIujwGHi3XRbjr2ZJO3jk3zMnWZTy1Yr6tVUSEcmi5FhL5oKy76MOkapEv
dG+KB/wf+OComei42yG82nzaqzo8SucTqtXN+xS+9np1LaqYSnyyg2AkFlXO7c1t
yJRHv55lCawEb8zHMg3IUkB40oAxbfz9Oo/stZtuv5avcFfd/uACf/F0LsHNHQ8S
2SEuA9Ysfy2yNrqsyQ0VauVXCNtz1K3RdiaJfMJ/mDSeGTHG1FzYAzpJcyuCKYOQ
ZVkADyXdQBkNRglYGvdGRYABMye16pfDJw6oLVuEzPX3gr6bwR0tx3hKbm9tDqch
T8eB9auqi4aLs8SknEAUI3lKNLRtBwYLLOh8Qtb82zJvfP5JKTyHnM3E6O8YHXTW
pff2WjK9P/fN78fDBhjAOZB2DwyfYYPwMTlIaZsGc2Hd/tXL7DgVh8g7ajygtxEu
mkwqzkrxNEkqz4NWgYRasQTViQLgir2gazuONqz5kPeoKKNIo4UJP83ZYQ2XzmjA
7Twpey+GpsgqxzmOq7fqOGJwCHk+uq8LCSrzXEhfADwqkyUQ/KmdWRq891WgbxIb
9VzPGLwayVn1ExfF8YZAKSSQY7ALKiSuwrFXHuJzdddbS+KSRIlopOgsz4Nx6SYw
c3/HrfAbiyYA9GP3wV2QbZgK7URtkIFzxhuWM3Mon2WDudKU1lnQZq6xo1WUSJGb
K01uLqRnhA3gwsYCZouAHo6p6WjR0DVBIml9jRFT1xBxTF//3SlIdAtIGfTvZFNq
Pjrt+8g/9AMAXNpp7SNkvEqq6r74tPhPXo6Uklg0Y5H5e6FqJ5Rj4VvRXOBbTrYy
qkrtliW5m6W62LEKGNydDTt0PRGnRBLAYWJ6f8Fn/YEGQjdos85s5FB/69dfAxGc
XX1R1SlcTu44JkThXVJWMHF4I/2y18ARI0R0UA2NMffpJvu6NuLNeV0sjYIrU42F
2NZDkXtfOjhnL4pwftyXGd7jWG//xUng9f4nxiQASPbeCXL37gPaHbtkW5gYHjzJ
7PM0OjFL5n/6Ese3fjZX4McCnElYGD/1FKVdUw8kg06WY6oWbUa191cxyfqvz69R
8YpVyxu9XIPGNwvCd0YTReYSSGj7vYhNMLA5ZeU9ZAQH4o+SoHkABzAuGj6GG99J
RZZkOxVVDh4nryByDdw3/LqtEY4F375LefbqQJX1UhzMaquX9hzvyepkfl4rkbsu
+KDAtl9lzaUrPnIvgRUPo5uw5Mi5Km2Th3kxqRjVQxlx9dYM3zPNF029SH8hVJ8f
h54J3rEU1ZUILZkASdINpO/gxD4tTGBQu8Bg8EhqT9u3NBykK2szUvfFou4284/3
3BjxEt176KZWY7hUEk6MYG+iETPdi7ZsuqOGmJs5WL3f8kAVlgCw+qcGt7jVKvRq
8rS2688jMJyc8fWoUFvhpZHH/tADq0zhGMPimFTcYrK+bxtJueSsuqoZ0WxC9qPw
A4UfX0qPp6c+/iWSfOSZ+qybmZXiqwFfm0JryiH4n6hX/saQMGbURuQAmXpnjgIz
ItE2jylKTRnfGPx5KzWQD6ckwt+aEZJzDWleL90GCFGmh9eWKqrb5n+zNssiHni2
CJ1W4JZUE9rzX78G1xZVVUXzl8dMGmPiyO3RmQ2RsssL2K1/j2rbEg0jiwAYjkGy
El7i9zk72t5iaqpATqacxGiZftqTVk1CS/xm3BxN9ebXimiBU3ihBQSGswM3W+JA
hCxVWhcSA6uQtqApNOGDoR7Ddl3p/7vNZ0+4q68sfi9fFsnrDnJLb7THSVdc+TbC
KbbxWLR1DEm1hNabcPZySVNJuaUIJbrOGKZIxgPzwoZ5mIU2foTLXeUhrY6oyJBd
3BVynXp7rOgoHTQwDZ/vwsB0ftrV6Nt9WwP/XSyV+iEMAQ5SmSHmCLyqvdNYCR1w
4RgsgB4/aLYSh/5qb4XZpr9bb1RIlLwx/BqQuGZOaL3yKDp1u1+IzbRqXOXeZIA0
0MAtezDS8oM+Xyr4uZmZ0O5nIcimQFiz5TGqg+3oHJ72zrEK31GS5ojnDg+dFrzC
mZ1IBY/Xb+uQ7fLGTQFCWDbO/hDzsxRpicqwPAUwZFMPYyjksk+CY0UHUuMQFpYi
4SV/UUpAJCU8w981av/st4/OIYlA/tkSPdBO+e7ro5RZIm8jzjqr3D9OgHeF6TGO
LUKhOVbbXOoJZaDgWDmXSNow0WXpN6dipOoWByhhbD5DUvL78mnCACA+7RLjE2np
vNf3TIXze1L/uGZWxbmYZojiLBhTIe9MpX33vrzlEqdUHAHyq5Zpus3wlTxiEbeu
OPnPA3RvWWMeZZKp0NgmlS7AO+cyYReC28u7bLVJBUOf0ZvGMkag5PNM0FvD/oN2
1CYQOmwE9MMhwSNsFtxUiYooCouzW6E7kB8JedUcZsFKp1Tg/7at6wsQRNUXHh7t
AcDi8/kPVs7Uf0UAJi+WH+HrvPRwlJ5icapjz2J53Fjd5YRyrzNEr2ipdrab4xGn
0zNPALlNFGyEAFw0tdBeEnixAHptPonQd4uooY5oxg7695VHnx+CxJ6h4zog2aUL
zNUi7KKu1SMvPLoHfKtJZ5Q92+VBcAfk/7SomphN5o9qN63NChVKRfftEnuK2Ijj
HCdqSKxftlbsFblp0tq3bls6G+uLklEXbKsm2XkE53pGv/FppK3xlY9SDWCJKQjQ
np/Ngku+OlFMB8rT8k/FAg/uPfUmcusd4XDYRBACVKqeINyoxPN29vLYjNHz9F41
VETLZIUxBvoHLz43VeAc0kTOvT6kGZv2FsY8rnFuYDJytPzZGEOYuMOrVMEw9XGQ
jpgV6MhG0rTLTE8YcXskfZmczNIgwSbVt7OFcDRc9UuyutbwFDm0J2B+/yYvGqQf
Smvx+PIpPD2AVw5ABDm7Efety9oWTQIL8uBPSG2NTiEjmAY1p9PKFO9Gq5o6ZJEA
D28X3J76+eesJBZwHagToNZkBLYwdeYpWvVRefZ4szig9ECgv7bcammM2sYLeW0M
JseZRG7+mfG2XiNBjgZRyz0vHu+WNBMf3STgbAQC300BYpplAcjILdvXQzYBmSbK
7iO+NLQFqYkSEgAPAWVgd0dXLA+FKcq+un6+QeOqbURTTO9eErrSKHeH3hNa1mzq
0Ao5t0LRsTu8rKWnKaE4Jo4gs9UC2QuI9ALnb5dmT4o+v7UgN0oDrCZizNNayiqf
ed5oVFhdl7yDcPvu0/O0YR6+LNMAhPZDvawSJ0rD1E8fETJJu39cH1Rrj6UfneM9
5w29Qk+bj7DO5nvS+HR+rtWo+ZaQf0u1T7lphkMObH51Druc0QUkRki6Th5Mrdhi
Whr0jWHC/CiLqzXsPHJeF7xWGlqTpJFO10xszdc8hiFNuAj+ihcvdFat2VDjSatH
Biep9M+ri/yVTZMufgcf6q85FnnRZVv2A9IoB3d1PKLbfDXE5fgirKu4nGZ7HK7v
R5u/pyBOERoJTSytCJkc5DvSBax9c96nV+3zPRSNddz6UARFtD6dnMoEBFcsGdV/
a24TN+Ua+cw4s+hS48NqbUpX3KoT0Z5tEEstRtqC8C3hHZ1ZQpQbfqD6IkUAbplI
R3i9WkpxQwpxNwZI5C/LfsRQOT64b1GP9r7fi8qdB2gfpouhdKsi+NwoIsnqNVrF
d4Yu6ePHQDZZissThJp9MUXNZiHQX/tOsYe2Mre/mYyASJ9bTAAJpLYtyEaQh8Bb
mZg4+rHNX3cGIXHRLbkrzDbssM02pIasP18LzAsskUeGQjXi7IWVDyqjEgqbGg7W
SkK0r+joemBsqx5EEnmJamwB9VDl3Yi4h7PnGo76LanEtKcgClk9GoppUGLWmiTT
etRJsBcTcodbYbyA/EcYUuJElAeX6dUKSSpzfISOotdRhov0db8OegS1fclbIq66
6LEX5YudkvHC5TSY6hx1+3sTLGwcbpfOKLwP77SV6XuJ/0wWhZJhZOmDkERQmnrE
GQJgMclt9FhzE8Zb+/wnPSQAK8NKVWppmQw6N9pHdc7RlZGNipwA9m+O7S7c4IMl
B38d8vX8ZH8n8g3wa7TTRlA3UCersrceF4gxj0HNxQZ1CDxfqByj64Fl5H8dIxH5
Z8sWZWBqRi1ROLyZ3/fK57APKC/Ff8UXfjin6pvTRGorFdhVJo8ekThi7qxFk9mD
sKpN8W9QOmbrji0Hcrhquszbfey3REr8/mxCkQgr+ntTMSNewRrS5fiWywv1Kyx5
RM8DIx9JcKpUcCU6QxEiCc3FKepfSBUqjtDTmveBS55C7UGczkkziHZLEDw4+cTT
oAnevetilbt0tk16dFrDBHUIonNghbchU0X6Hfbhz2alriWD5x/usKMGO42JOdRj
jvgC3pw/+N4At3bhJH8/hsKK4cRkRV5ImhRapDabs+xpK9LNooh4Qp6kJ7zu7252
Yro5yC14eLhahRNqgb4E+K/HL91VY3XvttflRkNwpEJDI6w/MHCq6kCaU4a3ICc9
A6cOxe2TKwdCnhcytK6Uz6SxvIp/lmgWuah3FWnJEW0DbGmiagdOMuoYm9dNaaDu
PmPZLZdO+Rjl+GEYQA9svCX+pY9PmtG+lSQGkK30NKzQvYDsAbL28ARe42zXZTBe
zYki9/md81os60OrzgaukGAoLgWNrB60T9P43GHfJnKj28+kmOL/uv40bCt4mnxR
UAmrqsPqhf0PdHcR1qVN3TDxIWW7T/+EAXOajog+t8dZoc81CiRvIlcoO2zjqkN8
5om1lmgrD3UhUptfEyOjHNY2+uZnb+R1TabAB3O8ggGwhQj1QX8ZMEvN3hDureAG
TLMwT6xZw9I3FY79KT6tjqmNXJxJz7lEwYmQ8pmjTdKK9QbNeOkSM7LcPGQ1lW/O
HMUHR2UNpzwsWptknE9aRXqz5CQAkZyL7O91aArLe6wWIexPYZPlNAkTc3JaS1jW
Gxme1PXW4dqUqLRF7vPW01cs4mKEW2AtTu9h3KR8OSbANR57HV3TWLW/H/IxiMjK
zgyWkydCOBnHZHTvdSW8/ACYAjrgqjTa/r6w3Mik5EI9mzb/SRHiRfyUKs6D/n6h
zJsqKEPxlixiMXOoAkYBAPUy9DigkiYM0OsdxVfahE4QNIs09+Gsgrb4XzHoCPM2
YHV12Q1Yz8BNKCLL9zUz4StHGhhdj3xTq9A/kPDveyuJK1u6DwSU9K9aq0Gy8I/g
3iPuXJYITtg7liHwOxU0MSnHQylEGG8UFNQVCmmveZOUTC+C2VFusG6ZCmRiYf80
3z6QxrA6Z9CcuTg3SFI2uXmBbVMUzn9ErGHvo6CWWmKrnFCZ6I8ik1Cz2GrIssgE
+AJAa+QQwsmRgEArMrW7+a06iSuEYD5gG/C/NoxSXPf3Ly78CDJ0m/sNg+VooihJ
r746ymvKEJCxbx8zMSuXtKrBf2OOB90odSABC25KXzv2j8KAXhAZmOT+8v2Kpp+G
9ftNh7cboTbx6yMDNPwsRPODhJTgNaX3Dt0CLDFqsV3I0tpLnGk5DuajS2DKcfT7
wIW7W4T9MS7i/YYFkxfJCNB4oGnRs3XZUHWxFyYGylvRr7Srbga6QdCLgyN+zXQk
ilhDGYqvgYsjXgs+j/p/F8ISy67WmNSThgaWYyKw6mOiiLgeMbsnEzLQL5yN9aVE
wzYZUzty7oGGz9806c8AKXaAjbNF8AkyUcsP9sEFJ6vflmgQl7KcDnTYKilew5OO
7LAZzjVZgkYRMuUzgtOfxpODvZIjQo9Sqt8fiyM5JBsyuCUW6PiNmQwcs/dDII97
k1IYutEgyJMPl1FX0B3r/oyi7ghqwECIC+eTiqR72v/FrnCuqRPGA9cAaBz/M4qi
kdNb+UypMuJ7W6598RQtqgjEnj8jDZn8onW/iz1HRLgqeAIf2F3KfaA9Oq/bkVi0
mrhWknyikoxjSIBnSnUjMJFfAsZkajP4/v8GXw0rtdgiTsszC+QuG17BMbVOyUbQ
QSwLpobsn8+raCWwNoplOmw8k8YzdSlR/09KP4HNMSHXGmNV8tA7SmRKaTh8Cqz6
b4P4VdNZHW51FqI6OnMXtRMpvf176oZ8x9Uz1JjWfB/6edDMk/A/jmmMi0zGnWAS
U3zE+KrXUVF1CCdV+4PM0XRmfhE/XgqaV3345vQoUfc6/xOnvzE/0D1Fu4SLQTJ0
tMfqFDuIN2luLl7g2fFz1/3aK6FxOKxeFUbYOEV8eR13SWx+mEdZHVgm1InLzP/X
r1ttFXsnMSDYhKKZ2VZNhiZPTuySGkd48wRMX95fPrS7jlAO6AuYS0Iy2Gn3wyUE
IqnADDIyQ9HEfKDr+ib8EloBBxTy8YixhNeY1LLwbqqPjSXKwWRKwv8sgXHvXx+j
G/2AOmakadCfU0nMzWi9kb9sNpvXJ7ud+SPbjNAUyqYOKH/HhUIZkb01/wPsJnFh
+IV+XGaiNYZEMwYU2BtWvdflp+f/tFcp226s3eygyLGxodhpKFM3TqYep2XMP2Du
JR32Uda0Ke5dx08sG6862kEa3GM6WA+gN7yEdJJEp6LbknbpRjwgc77NrxnJQA23
g5hbJ+JREtozfOycF4O7xCK9Y4Xw8K5hXCi9lM6J/f98N2eqLEEQiTXHRCHb6x7u
sKdLmVNBrgz/ySQ5x6+z+pBnfvSu+OK+etH3f7b4k0k3gkZNXBZ7jFLLWIOBdBQN
H0EEwp6LcUU8AQoyu0f9cOLkB63oDxcMwKa4XMwp5yy51YCSyagxX7mOE1csQvVl
2C79RGXWZhEnDolFqwlGKX63OKWN6Gkwpq7TNhhyrEWdIcWyB2YRvRoLwPKpppPa
6D/yhJ7xSHf1pwiS1jb+5ZCyndFuRfX2P+VVtOCg5k1J4T0RcncGVX1vdXlu6R25
aUCH7mmyC22QxtWlOv1oZe/7SvS9IOiOKw+nZiguHqAxc8aA+KrjPKcd6gaqXa+f
G0FjIE9aZbq63h59qTETRoamCui3VMCpK/GTU4AwaEqBL4g4nVE2yhospRKuC/ko
XLZ2vNA2qjguHEKoy3+QVw6kEh/+symXTae8dSuiPZ1bjbIp/LjaEqQOgGUATepz
//Ajul6SODjr0SHP4VnyrW7coSkjRBVKaVIAli3i64Qspc/nrDYb33dELigU4yVK
VLEAn2X7JET78QcN8wIK5GO+q9wtPxKZxbcjdiMNgoFUEIvft4+nGY561nSZtXIL
vtY3qn2zIKVT/PYHz8zirWpNKCrmS3PqS4UeTCvKTJAbM9DZ/xVP6CH72hYl0zss
rOo8bsyL1CLdYvRHjfhVPKvOc7+5JAa29yRdMKGPMvN0Q+tehEa6UGYuW3F/6hLS
Y4Jwh6Y8px1hMt0B7bn1MISGytZCAPXJXKucLK5b04+8dNXKbcx/T5Wvt7iXO3/Z
+TVWzqBMUJAXoTgn6hoRR0dzAoZvK5Nfh7/iVwfvGnml3ydwBLi7HYpOZfoqPwX3
5I7HWxq665Cv6A3uUNoe760kPD2xFMhBeY+68XzntWliut7USi5qhm6x5upWrfb6
9a3hm1YHfVGsata3t5flU0xpDJCy0CsIhB57gJqUMpDi7G7xGE5b1Hv9uzAAma1G
mgp3E++jmb5runUu2X7eokqoTb8kvOGFKW+d/y//u2vgT08GsVNvK31zwpeu6rge
Dh/GRXdzoEc+iMvEuAbPIZu7SZ8RQm5rwfgYLd7+AvhHzSDSrUNRVVjso0LHSy57
6p5Nj36CNY45O2xo4xQZBy4xcFysrNv5NgcvSw8aQvVTR4pXG+cpr89ZynG53sDX
oqdCRaRovxHv7KgvVTCbtqfUjWgURj/82tI8HHnNmfM9mnn3+Xk6PSZ5Mz3Py6GM
bOdOLxqcZpyWXbhotXRSJGc4+rEPrp765FLPci4S+FpU+8PedebGW2ThTv5R31p5
2lArtVLbesQBbADPZvEcPL1ulDpoHy5wY5Hyz7z4W0bEedlrHMcb3ulPD8Ephd8e
iv/P2z/C7UGssAxiwFjSibV3VfP6fdbeq4VTYyHEohALdzL1+8AZ/k8kpg3+iKGQ
5fGIt+rFHEl2oULLIcj6vlh9Q+q4rKOLQjYMP0w5YMzlT6yQEFtShz8i8tOk5+Vs
fID9Eo1OdkeofcHCH6+rYp4L6LyW4HE2D+N6OoLqTZOIclbjOdNTA/BYtQRLxOv8
tYWy/THmFCbPyxxlgfjsdt5WSp5gJ4YIwdP9btc3jczfQoszxPDqjwL1fe08wrXw
bfROjtKmhEh8pPqdjgg2cM87VSVauftuqiVdH+tCeYZ0YY64n9XAaXgOF9ThEnla
tLToqG2fTh1l/L3EGst4D5D/faktfP2uvAcDBkqXCl3Ys++mTx1aoLtQnbvncpM+
8yUwRpfdbgNJkBLnIa+2q7N31pCHUk3ClqqpIuf+z4aQLM5p0lPXxsI6BqQ+ikaS
y69Uu/hgwo+l9sU34pICt8PMM5ObO9NjW/pMSPfYqieVPp6xTtm9iEeTR2M9RJg5
QxbXd1bK+xO0P5tjUbBIsGBax2vPv1cYQ7lQPEuJGYJ3kB3Wc7OXz7tyihAr2UzY
8DTos6l+XJMxnvp6ksx5PKf9rDPEeoFCU1kczsKkoZ9FW7hSVTGkoSI7sa2SUG9M
gn91yLGJ2vV4hnfhR93QP3eCwr9/J6/+GB+LNog/vADhgjGuop0OkDmdFJV2UYu6
CsQye6o/ONMgJlWlkGWc4TsIyab7TgstG2rbOUmBFmGUMTqJzt8ynfhSL2Myqa7g
JueLA/LHDf0n+TSk0jkBfkr5QIQwSiOZGFW0Rcf5pquItGT8u038MEcg7EKSGJ+b
thIFg2dB00errOQ2CTE4Ve996lZN5vJucq09aMqmsUrsuvZi80uT30If2/JNHbhL
VLx/d1ya4yNGbkyweHUp40IXf+VLmIV2fBiGWzyaMJQ3xX1HTFLbLc9SpyTJkGRH
ffadmYsByGueWNo33W4NsqnWMpMaZXnMzxKbAQe0D/NGg9dRPl8z/itBU33qXa5L
JR/5BhpFCYzZpJ7xleFBT+cszQDTNC933gympiFTnBJI/yE+BVZ1OHyoAmX5wclO
/+mSUF3SiAFnXKMMPGhX3f5V2b9CsuF+VjT0j4Kjxd5ai6zwm/3DydC+0WDdC1Z4
Pny3wcYEwOB3bjYtLNtGdE0g6jMNzOImti5EdeEKvUh+LTOx9DefIbbgAydT+97q
6kIn/jKPkZ4xQrLVn7vasfLKaDzZ+ka6sjCrod7hnzydLwtPcMNUufRHX7GUPWGr
Cs/AJoYAtqmVAPwkghH8OCPmjJLPvpGodwm9+w5srZUNThY0eLtPpjo7QvFO4Mg/
t+Ns0lhS3cfA4isF20mgYUCuPE13Nixw4xHoC/2F7/zJ6m3UQVblXevMAr7DNqR5
7CyAZnBebOhlgVopWuACOYRQeMWfHxJthLozKazM3buBYJOywD8FoQyiuOqgYHql
IGYhPpNoIRB5/KOkOYTpHJbFvuZlbbEygQmB2c6Q5NJBFOt4vI9vvZ/DtGapOADc
48zOtpgzhhSiQN9TXrf5YZgO8XluE8fZSvMa7KhSUORxANMKNVM7DJZKt59020d/
mzq9PXOp0DMY6AZO85etoEt6wT7XSaDyOhs1MPddZ7Dp0lSTS+i9KEcowlApSsnh
fVZNMRVbmegpsjTai9Aiuxod5ySxL+2XFI3QkgUXmNj1IgjfdttLZHJyEnPKihqD
QlY8jejfxSmMCJfGASx7yzKxj1fICJreOpml7ehLTvtyDSA3yhVpzJxz29hZePjj
V0RnssbTLL7nydq+VffRcouRfUtErDXSsuDdjZPuXZLsQOymxu4X/hddg3YBFtqP
0eRNjctHO/HxbH72dgWom26Zat+asJjcOzBoWBb+k8Og93gfC5Gl/Zp6L3zgVbuY
KaYABaRGex9mRDEBfcUQtmk4cB7DpKUfPlQkEGJn4BRS+LBQjz7ztoSJZ2v5T6zv
3o4Vmu6DbhSeG/X3gBa1d+0IX8+85Nfd4P0HU5Il1SGXSrl78oc67Xbbiwq2D+ew
8iQMx7Nkj6PKE/Yr8O35bwtcsYh8QnnYjoaRwa3kCfPkLPidGu1ya9BWks/VAmiv
PGp0X9bvLSJ4KcSKvNcS9nVKie1h2m6g08fnSHo6gabWswFuXyHZiraTNJ09Z211
qo3+B8ib51xbMXYFypu64JU1TmfpWlQPo2kHcKIyFWFB1i84vieWgvlLmPSGBzop
12RBjvfLYTqSHAF07IWmlYmtZ+sdj5A1ch0tR3h5L62yzp0xW/gt33utjixuH7ZL
WkTIdzqBc5M8O6Q76393Or0YTZYeu6ur6VmXcwDVWQ+zbvRk9sqW6GCy5gCOAxcO
/nOkM/7d8SY8D11/vrTBGG07rZ4C2XUoER4pfPIL3kFqiK4kEL2C/TxLMz8UpbMR
Om+qyz9upqV4ihKgeuJ8FHr0PycQXHwGADtlUwsTXBfKddLklxMOzfEuIIAptsgJ
qcy8pOx37HHHjt2MBHjPnv9TiHU8/uq2sJkHvuTXJBy5+DH02gveNKwbr3Zm9w1A
tiG3Ik6L/mieSdPBiem40K84gAqsM3r2rrhacVfeGcjOPBRjG99H/y2pNbKTMXGH
CFwywEo815T6eDEa09tQwW7+bpcwBHMGor3CKZdEEsJATd2Tt5PKP8IIoFHQENmK
upCbKok4yWYoarCxG8QM3qJFk36GCqKV72CbvxyRf767wDyefUhqsR8GFO9PDF3B
S56sYW+9u0+e/FNk7yD8T89FuJg49WX3dZMQZ6JCMJeFN7EHq9JZ52tzBXd0Sza7
QffcYXQ6ooMkrzFwNVCuCeepGfbBHznjvRquLyZEbiAGavAH3JQRh5VCHgQy5cHB
+JA9ieRaFWEg1BpW5l4maZpjdnmiYqDKU8S/jKE4HdXgicwwB23NQZV1DdlF5ewQ
6FC2EPyLAzjWDKfFoyIWwhtaKDsvQdPTZL+hoZcqNAsDsGXQ8xpYjEeGw8yHddBt
f1l+HJWBYgGxujkm5pSk8ZGn4QMkIMSOy9SaHH3Xsjos5FgpDF4MVbURHDmY7wyG
v0PP3797q0K/gwpsPADlc7HZH90kPJKMU2XAWd/p8QCAUbHrsdntRNxQFRcqK305
CPEvyfVN0TKrI6r4GlNKfeikThnSh60rkGNt7n7TPR7e0O/0PjiQVttLM+gOQrUy
T1nlH3AnkJyRR/hxKNFOZ+5bVz5zyeFkLwG4WgVObXQIJqD97WkpkRLetFrbncG+
Wspb9eP4fJQJxRvlI0oJf0N0JsDh0ZGj0l0uybO42KI7iBKiOR9pRk9W4huYGEOY
/NJgWQUz5/l6RQgRAWEzTeSIo6ut0cF3JejlxAbbVll05op+DMLgFx1n7HpXUgvl
A+saw5dTB1JRKTxNAsEPfHAo08Ufgikvq0gUovJA54KTebKPGnhmJ2bfw7Oo94uh
RxPIZ7alE3Zi/VmwveOVKc8d233DpmVlnVhI5BPcvg5TqtY5wuqQILI9+H8M4ki1
Pr+kOiZAH7Qby2w+1HgDitdRVL3cKEq1nWc3K79PuFnEN69OV9LWXVc31h2m1Axy
m+UoIsQJQPWzs4fliotjVO/k4Yz9cce6VguHcI/iDdHOJXd7iB9cyoG7vtcKEURF
YqZOh8KhGZa/nDhkf2g5tdxm8XOG5exEL1tdvH04zOSqixOaG1t6DB6pP5XWdP8s
GLkG53q4s98O7oDlh+JOJK6YgoPWdl1dxVY+moYdv8eLj+n2zzysxEzVKdVpY9lv
U4bjgj/YEu+qgBOE20woBhzq5dbzehRNfPSRirIZKyVE681KXcgXy/7AlHStzb8d
uYzI8OOYvL3ByoEgEmXwigojMp/tlqad5cynHQWj93Eq5GuG1FwX1V0918iI3VOL
iU68+TFzXRpYbImuph8RK/jM0vWT+qSdiMOtixAdg117vOnfiG44as5HxPiN/b76
5Jdh/xTOhJjJp4/dBnqPWvuzCCOs0lTkYf1gXObVy7rf2EkR/Cdwyx6rUf2ld6e+
eUfC7mayX1osbWbHCpejynP2VQ0rlADeN+E5+BfRkrxmnxGcYeghhC+66Y50bnOu
IeG68PYYeCMUO/neerpKeBRPPDoj5ScvGWVHRFCe/UekT0x1r6eAAU3jlYHYJepN
qFvQ2yyd7i7EK7ZJWzbp7h7xt3aXc239mT2RVk2lv30C4sfi19zECaS8zVyNaWIT
WvVVmgEFbaY4wUYs+81C7Or+LI89UJZFmpUfFZRZT0OcqxKGjT+TQWwiVULnfaL5
w+2qeoEz/LZrJSnNOzt4oyV6Wb5PaOKYFmBaPhZsW8DvAHE75IzrR4ozeyZZI6yA
ZX6oTe6TAFOb+6G2obzEu3h0Vy2AJe9URNmv7l7IkUL9ZUXPMb1gB5OOReRW+CAv
vzWN37xgUZAnuYMfTe+WQMgC513oaclPvdEkdHx9PAZbbLiIqpXCSHZjw6T9uOFQ
6g/r2IetXBA2xqqDp8ow1wGusksN47lmbLJdWNJT2GNx2czlXFCcWe1oLZ4nJf6U
sZvGoNAfg9oXjcAdA9d+z+AT/X5Q82Ob8jeipDepl9jSWJ5qoe9En7G6Fi7TrMvN
N06FrqQd9ZpU/BvCKtHcSu9PWOhs8I32yJDNO+rn3zj3a7YIeppDYyN6Lo3b/hEB
9SX4HBZ82BCbPOVHnVwloQxLBer5ysoQTpA9+L9Ldz7KEzg1Dgj8ux3r4sLKsxF2
j9H+leP/jBFhUob0iNJxliImpYx1L+B+PcodKL/Ky9tsZ0stYWaL9MulMtAbEMwb
tCZZ0c5Gm/c9+cHiOrTiqkM0Lk3sT79hIJhNQpeVwa5sHt16wdYl7qgKDK+D/ctr
2aeidkkCqjyUQ8fDUqO7Z5WwxDSwMEeL5aHZIrLTNsxex8KpGcw1mgz6UnwjW517
rLe9QAsDaaU9NdDZ5HuigEUPfwSV/oKC2F+JYxnEFJqmstsZDVNfWWpb9wCy5k10
N9++NdUCImCxAYll+QuQAMYVjKy2n+8t23tr8ESeSaOBEvS87MBWzO+3CLbIStX9
vqbCUgDHtZzruVIwhcGtrK5QyPpL+yj4ubUc+izTTIsnqNTn5HI5aO4JN1+M1ywg
`pragma protect end_protected
