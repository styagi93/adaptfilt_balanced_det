��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,G�ss>ʂ�C��S��D/��mD��J���Y(�H���U��B��Z���qw0�Kǿ�(�yvE�e���>�)���L͠^����������8�4f.�`9�j8�.��ٺ�>�q��Ju�sUE�2�<4K��1Fgݬ�YxMI|+f~�?�Ԁ�;.msO0
��*OZF��0Ǽ�|#2�tц-bٶ���8fJ`^��U�B�$��~�(� a���xKX�!�u�m�T|�"���M6��zf�q��� �q�+$�Y4�����A#�u�.0�*�",zb�ԭQ$> ����1�h�XG1�T��w�Ԝ�����lȣ,�J�)u0Yy��U,��󟒊�<�<��m"��zA�˲y%���u���Z[��<���s=.�ƦkC�|�@Cq�)aR���-�C�-ߋ�W�-�n�C��������U���ޙ,	�&�:�Z�q"v}\�J��lR!^w�C���UC�ۥ�qz�C���a��u�)N��}6�o��AZ;�e��@��D���'��ZY�\-�V�䙅�ʳ��Vw��0���X��aI��W b��E�aoׄ
����Y�� (���&D1�À����Z���j�Bwb�XQ���j�yAE��ul.��m��R*L�<�X�8�T\�Y�,)��s�ٍk�e��'�)��M���I���{@[�͈sw��<R4D�ui԰�wpu��a�A�\]��N�su������qCQ��,G^Ӥݦ���z�������2r�K�SȰ�DUE@�Ys�\Ohk.9l�͂o�ʱq� �y_���G�� =�r�0[���ژ\�C����ӭH��3R�	fA������;�� 7)�}&<�@�w�u�߫nC�)�3Š����:I�^�U6�� �i�����/�W6�T�m1K*#�P�+y��r��"t{!zQ}�	�j����4�US7�T�5N��7Rع��Nb��D�K�{s���_��Cٿ�H��e`X���}��.��8�#�+�{n`l���#�����Jh�	q!��&�w�e؉;�0�$he�Kҵ���ω�˺ɚ� N�ee�boN<p;�s�8ڎ4�S[�I�)^7U1I�`E����k�x��r厰i�� px��d�
��u��W� S������ģ�=�d����B�\T�{��CU��^�R�Ze��B$Tŝ�ĵ0��(ׄL�6���Q��cg�K�P�Zſ��l����n"�R�M�d`V�P�����@�6��&fŁ������bJ�P�~���t�v�ʀ��f�c�PrK�yO��1�މ�L'Sg� �,ǖ�0�!��p>xk�%�q
jB-���V �ɲ�}YEҙ��D����:����OܕEo×�!B�"�4W��A*B?�0V>�;����:�f�����X߹�b�_�q�J�+�~T/ �F��b�ݳyl��6��v�����a������������l���x��)�d�����)ዦ�0���fw���ȗtD]�t���0��dSYi]S�B�֩�i�ǳ�kIm��RK���6��!�g������:����p������X��ࠉ�x��qu��U7�4J�8��aA�`B�2f�@��̯<ze��y!��v8��.�Q����{16L�HwT����W�)�4eJ!z�	����N8�H~3�Y�O�����F:ʓ�ȶ�jDĪ�~i�{L���RV����d����\(O�d�f���
�_aӞ�[%d**��A�wj�s9�m�!�>��D����Qٮ��#2kΛ%>���AG�r�bk��7����pK,�ۍ�BY��3p���{=@����g���)Dz���XΉ�qu�Ωo��]bA��ό�haƓ����]��A�O�@��4-�KP�M�&�^��0�\�@�I���YtnJb�b$t���>����)lxS�@t��U��|�%�n�-2�?Z�i{D��G�i�P ��>%���ߗ�����O ��]����L=+>�S!�iI�2D{����2�gF-�Ψk�cx��+�<�U��-�H]{�j�(8�s�3[B���9D|b��y�.#/Tru˗�ȥ��m,7��a��{�y�TFw��L�a�l}zZ�]:��R_�l�v�'݄��/^��������z���t��}Z�Af6/�N*o��N�C�q��j��y"�R��|=zV��V�8���ۚy�~��s����l����>�~l�0BA
SC<�ʛ$���V��?&nH	���}�s½�{������;t[8��pm� S�1�dNZ�Qz��<����U�|Ǩ��������w<y��DPRDa��j!	L���a���)�<J��X�*�s[����֟��h�쌞+�DY^���Qy��X��0y?�4bay���ˎ��ST�Y��j٦%R#�x�x���q�/4á[�/�@�����8 �9��.m"����o/WP�j>���u,)o��|%mt�@�!(�(_�n��W9�(�FcLU_��/�#�X4�Z�R�հ��  ƫE����r2��UNlW1�}TH���t���ye��m����A����G���u��&>6K��Mk+"<�	D~�@�C@8��(�t̒P�M�\�g�2Â�.ԥF�oo<5J"^	5~+�����Գ�v�{ ���Hc�
���3���4��^@�cԘ�S��(�{���}�gT��s!��hx��:��z�j��=>Nai��>�6Y�b����2�$��Q�u��R��� �Hڷ	#����w��'�2Z\�:���$��<=�����dq�w������]d/���N��Jz�P?6����D�%������|�'�N�7���q,�����g�:�K�ēI��'�*0%�29�JB����Z������[�r����v�yГ��a%��5���o��Hi P�?����V�v�M�Af���v�͜�:���D�4���58J�:T컡��{��#����ۀ�ű��',��ߪ�f�G����r�Q1z*\8컆I|�b�p�K��G�xk u�A�F�W�	9k��E��S>&���˧松I@��HC���6z+����}�<|���K=\IM�^Ue�B��YDM[��.k�	x'��K����.v�ox:�R�v�"��L-�;;�P�*|�f_^>J�� �zw� �JjW7ȥ'.�c�m�\��
(�P"��d������^�;�o�\�����f\�N:��aW��1h�\��#Hý���?H�j�i����!rocjc&�^�j3_v���$����~C�q+�5�,��3���~%ˡ�9�ǫK��9 ����qD�Hq,���[4�g�JKhM���rc=���,�{b���FW��lkL��2�� +:f/7�gʉ��Xx�&�l�a�k�i�00AJY��b_���/Ly\}+���x g�E�G���2���\��D,0[MŘ����^��47�P���n�K<�Pp�q���m�rA!׍�h�&@Z땆��=���!?�T�１��<ң�	��3�p�����%x��`��6{�ƿ�m��Z8���
e/�JU�'n�P?��އ�x ,��� 8�q��|z�P��5\&��x?ye�q�h ��a�+�
Z�n��_mk�*�L�%$A�Z.��v�C�V�� _b���SZ���8��Q������4UEd$���RDZ�������# �_Yu�{��F�}1���8��˲��a��ü6x�����;� ����:�y�/��,�"�>\']+��tr�-�J(ΰPz����k��w�3����얎�(7A��=�շ&�AU��
`$����s��Ѹ��[4�B�6����x܈_��
��ǖ#}@�)q��_1����'_6/:���E�t�H��'�r�hz��cAx0�*���y�;t;o^�z���SJRL��V�9ULd}*�L�p�@�J�,�˖����&Y8�aܽ��i�z��A`�#G����쨲~�H����|}|��đӺ�l�.:��l8����8�e��ͼ�����C���릍D�kp��դ�{2^[7ɶ,�(����w����dvd�y��,]Z)�Q�oo�i��s�!ći=z���4�/XQ9-�4c��O�rxeuĦ���]we �IӾ���޿�0��`�p�K��Qm��="�i�JPK��{��o������*&�GJ-4�(O����N��Ǻ���m����n:��Q�JanA��ڒͥM6����ҳ����Hx��A򑩖�H��/���QSҿ�*t��qe�:�zd97���;��w�w#7��|�/��8�W?���3쮫_m.��{�����^#h+�St���7ߓm�����-��=�)�ą~�6�`��5վ匏[K���;9^Z��M�W�ـq2�����������f垀^���V��ϗ��`����6s��^ܽ=�ۚ��?H�Q?Fr���-��X^�d���w�ž�)B3� �_9��Q�GB"k�Ҍm0ҭܭx��e�zwaa�m��u��- �	-	��R�`J�����2�0�a�ťq	vqv��])oDLOB� �U:��jtVz�:(�M8���@��]͙I'D�8Z�)�*��,�?�\����p3j�⟐�H�J]L�Jm�6��i��0��x�4�F�~�H� <i���htZ�ܽ��A�l�ԑ�%s�ߓWћ�2l9c���r�:���:��i����2pN f�<M_���]�M&X+ȝm⺨Û�n�kR�c�ճ*��~^r�����"�D-�+s��{ۈ�f������K�3C�A��_9Z�(sT�% �����q�� 2h/����!�=��V;mT�g�A$#�_� V"M>�~u�"�X1!�b0V����{�%I~�vK�#n��e�t��١�mII<�1�a(��_�����I�u��|�uv�W-a�~�I����e���f��a���a32q�w:�W9Os%:�\b&jl�:����MD�pg�W�Cl�s|�J�'�����"���;Slf�#�T�����*m� AV�ĩH��H��W��)��鍌��N���ޛ�
c�9߽Y*�a9���7����-������zݔ_?:���Z�= 9//v+���XpاR#^�����]$K"����r���r���un1'� ����R��ih{��Sq���*�
�����5)W+z��g�H���ē�ņ�r7��Ku�G��C(�$�C��R^�=!3�pHH������ى^�k�`?��)W"`���-q�k2A{l��*�HH���������p�"7Lil���o�� ��|����)�٠|Q�����.���P��������f��@G5�14~�z�5?��ߚ�����D�I����jU�qT��KSk�h�2�>��Ԡ����Kw��.���^,>b�^���gdq�o�L�^`���o��e���	=vJU��$0}E���`�/{�)D���*�]�o��(�ْ�e�'egBvݸ	��A����/RK�P���Z�K�D%��x�8-���)�z8�l�����Q|="!�yC����tʄK�y�t��I	���ջj��$|�h���h��4�A�Nu�uG't���$���������߅��2`}���WD�G�h\���7��x���>t��XY>�h6Q�M&ŘuQ������Q
����께,q~��J�7b�X^�(��1p"�^��(��_��  �LpL����no��S� ��}8��4���n/%^o�Z���(�he|K�� ��Í@҅��ӆIQ���ɔ'���?,�A���$�g$�:���U�ٺ('���|�_$oo��q\��֚����%�4������]}�/8�y�]1�'�L=�uA2�