// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mjQCggay1VH0q6ujsLYB1Lv3m6DVPORk2n+sMo1jjfi1WCn74bZSI/UJzM4b2WR9
FvP4aBi2nCd+JRgGd7IX5zXkiSouUfwCaKPdeyoaLscZsREhB4fefgcLAHbHtiGQ
0VI/I51VsN8upOZPA929E0Cvm8EANfNa8jhAXKb7duY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14096)
1qywG7zll+6zLs9SJtRMFrmkOlhao0swZwPXSL6ATaOKjTPAVd2NZIFLdOAKgq2A
SjEx8qfACk5q3lRDh+IhVHagLfvP6gNqTRW9N2a5F/94hdQF8U4ynSLtznqhEuXm
bkj/3x+4Up5isErR9Fc49hWQAFRmcdLv6D+iYphRWRfBQJmHNHOCsCjxBK/Jq4WH
OJV6XhNP9t34R4OMOPksgUdYIgncCo5ywSeShv29gNi8fgXnVwunmXf4ZnqQM3ZP
UsGAIY3HZqhukNaPdgrgt4O8p9PrwwaPsjeJmOzwMVnrnro/IIegeSyXQQ5N51ZC
/aEvMnKVeyLpN+s3xbDD7iI267kOzijYKgEFuBksDZUrMbt0XZKTX39rlEhwVkYN
mZM6qFLQhIVXFpykFbSricI0NNtpIDOw5br1m+I9N7X7/jBPOjr7sTXt5m5sy0fN
/Rt85QR7q8Cx/32VEBCbDrbVj5Pvjpg31uuZoQJZaqiytZZze0j+mdIfBVXoA1Ss
BXcTV70F5IxrulNuzvZ3ekeI+GynwEh9JdRrWWW/SMhbVXOwobJJsKmmshkpDrQz
6zBlVc7Q6aSTCG+nibV9K5OnolOdKrvmiRFWeLcbzD/sm5CtUMZ5hB8JZVVlpPTI
nICPs3S7i53TAqNLSEUtNsdaP76VfNpvTXKDmbPQTXl2f17T2lJTXK+ZCTz/H1T7
Bq4nywDqlAAOBs0FfSa+TNoDdCV67/dWKDnK1y39YI6A4XWuAkY6IKp8xgqc7qQf
Y36AlpfeLRuSPrdFxKaxEHWh0Dx1K57A4eF6sh0O5JDzYT8jh2hXRzCvw1800K/c
UG+IQMgL3VqG2UBas6LfuxBF6ONgN54oVUrv0jUK7qKlvRg7r9J1g0tLWAcANEIn
YqZookudiX+PLA8EQncp49XxGRIj72Unxfp8Mj+pZRUdLEh73zrUrwvvGbiFjQMw
IpJYu2o0ScISgATVcrhOZDeSpD+Lk1SOsVDSP9JY/o8gyRMN5SbbJwhm223+7cjF
acv8IerFtXE+CQrmUeEV+pSQxy2qOnVeRV1oV0TdZUm77FuOPSQ3jKMKhw1QtvjX
gSpUCiiuoqIRCLXkY8jQG1BjPehneJwZ45+MR9/FkMFccjfuncTWKxZy6zvKkfc6
CK7Jefjl9B85m8IsT8kbGFXwMuk1Hp9elhRQ/o9APQ6WFGe8HXMg3TCMWUoPtHVe
ilA5TpyWMpb63xBTKE4CaesYIFnGiok4nvxnHqwLOAtXiIH8oTohM7XINBeX6rn0
89byvtP5Y1ejsTT/PucplDsdN/rVN9q0IbjhalN+8H2YXgq/geJAYl7X0qNJPRt3
g28dOFYSIr1wHkQPxGJ+DgdysHx1H2Kn+ptncyG+qpknO0/MfRDFxdp9sbWbZTIj
VNrPfHTyoO3iELA9Volft1X4NcAGDeFsgvPN32CYtYoPS5pMIzatMXYQpVrFL2RO
VwGgEGiajOVH+7Jh37sX8tJmG+MTqc17A1NLWM4FVoUf5HKKoj8EaI7Uin0GP1GY
MxBtiAgb4z8fB3jhQmxYV0+YT+R38QwT+9yKmNUkbWG1og3hR4Gui/9fQNoNMYUo
6zGxGGPfyZzlAlOvMOrIGoGrUPZcLSVzkggNoJPDVOmdoeJAltKfTZ+4vMAPnP5f
t+8CaqoYTE7XTa1saNwnuKhImqhrM6g2nh3sJOkOpITjjEF8fdgoN+D/mJezWjwg
6uRftIMyeHJnpJfKv59u7Xplm1/GZbu1SkRFgSEYVBprb6G2EA37KkVDQhe9B3cq
9AR1jyjsYf+ZHsyK2HfFmZlWFHRg7aCbqVvkQxc355OBdwRXWUhrsZRL1lkLWF8S
5LmEY+OKPDUuyq7A0lRNs8vdwRz5d4xVbnaCtXbzKZMiAWlOjy8fiyXdrCQfwW2A
W3MLNwNOwwRHuIg6qd0bBRseuxZrdL01NhKvIu2bT2l7cp2WYOoMt8aravNE/NzK
7udY7dJJ/5x22LUfBBR5454DGXFobgx+zSqT/CPGCnYJ85uwJebISRlKdut52Ca7
1zZWZFgYiJ3PnZpCb9HE21coW/yFLdkM23BBUfxthG8c0iwAGtJQln3MNirm9COY
0z/gVdkzI9dz1doDMVHvM/z/MxBhEm4XdTU3YGKbJZiCNt0QKiFs2s9XWhyTLmq/
h/e2IWIDHmgCqTZM2O5hYW3x0WcQYam8MyGSiaiKRuQ4oF9q4SokguwhCIPZo7+H
SfV8iGCmfGJwur6qF8Ncv66MeEDVUZAWH1f1rU9tZ19RHLwh3Q4DqIEf1YK1Uxon
DSDq8ueOqPojTl9257oXAySj4nnFIV1vOQpWGZH4Vbdh7L282ExcGylDOyC5BOse
S65aI5oD4rULOBWxCWkrfFsoGo18az+tEk6DW4hwkzWAo9TuDrkSvRZvlLY4y+nC
THIcYs8Lku9T6cfsxPENyHy7AkXGt6QlmLlzrEs4ryalKvCcizqAoCClU4q2kapC
fwrKEgljFWD7vRc1J0KRffSRkFXdfYf7nKnQ2nF+YBtwQe6J1HDR3J4KFFWg7tzI
xY1nQ20WS9Y8KsrzbdyvQypOGVnFYMm5UUhOcoZRBfCF+t52eA4R1NzojX4LkmWW
E3qw3CI1skwvgFd/pIS4VC55TND36NDScXtzF3MLnG5aVGisY4bQADp3+A7kCIb8
TTUDw6M28jsEAYd8QZHzZiIVInSv7TC9XhRugzbtWcnMywUPSf7BGgoMf4NkMXBr
uxcFrOw2qtjub+gef+5pn8zPjfiwRZKA4JsbsNgHJn25yJSERBeQFSXUzGUic5jd
YEBorYBnwK4h7/u3ITUyKxPVdglYoIC4HDV0jNEg4yfWVBmrAbgVrgJrYlbXJAdf
lJeaVGFaoIweIa2HJrIkLTVB3TH8cbCVipFsXii3NsoUmtFugTJBmP2lOuY0eCGq
VCrSrg1bBuYKaZ0d/CKEJNX9dTJ73Q/jiI1QD0P+jTRjUCfMYLIcykaoKx0A4PYZ
Nn6mRhxzix0vu+RvY5aahXF10ohMbvaxmrJHufyXONwfDda38oGlCnkh6VSkpJpk
zGz5yScmMPsCSs20D+hkFi1baqCE2oBjYfVRmbmUTdDXPL6d2KWwj2qk+OQHmhe1
ZKm4Wi9MQFOBHDhHJ982Xvg739RNd8dS6OSe2pWXE2JrfwjvMjcNnOvKw9OBnHYt
XbT1yK1hckUFOAkyWIMMkS6uI0ursZkaLMHl7lONf0Lm0PG8GjihftrITJENZkQq
uV/RHLj/Vg0irdLAsC3zTAPH6r4N3pdkMkBd7C3Sqfxw0XjKMs2JEsz2ASbRMEU3
xhFPPUQnem91mw/wB0qN84kBjMikOfezYUd+zV/8wCMs7cWhCrAGMw79vZkRjZid
WxuInztNrtVv3y8YJB637zVqpUls6zfaVRRowv2q5l8sHw8aiyQBAtbj1hBHpUsO
tlGehYKXmCdGiMHKIC6UV81Aj3sDjG1N4YTVlUmR5m+fjCQr0nZ6KqVFBmElDWRD
oJYBb09zW7yWtq8IQ/e4ffEQEauhhyYlEUR10uG3PZ64tt4syRSDAcVf6aZpzA4Y
ObZv0C99+mCyhN34Yu4mWLSGvWnqFBdKG1a3b/OOlqCA7gXRx+Gk6/D2LH2kcCT4
Ry1NJROIRE2vyfHnvIsbn6xDmFbd5ysIwhZl5WViiGQtUGepR+wpOZn4n1U877cG
RZ/vDc9DBH8ajgx9301dc4z3yUO6fj19uGEwRo29aqq8o/bY46w+pfk/EcOZaXy8
iw64fgYDNoZWCU2W9fhDmr1co3X4uEN3y7A0jcLYNTValUJFRXnm9sN9qfROwb8k
kDE1bkVD4WGf5FPZZKD/mDg5j4W1SO7MVOAi/rgJuMq88PVzyVKIlmedbnJkXZxQ
Q3Ap4OYj7/Cmz5e5Hx6IxCbvVpavHpDuW490jVAyW8YXcrTXFt5Lisn2Es7XcSE/
KYD5QktZ7VMLKF+nZtHyZEJQOIAcMXmjfKo/HKAZ8hjyuIIedecJGn0ug+FWndmF
n4JMyhrtu0hGqJ3D0zDy34VDUyu8K8XZjveBcyFd5loHt/3wKQ/cYlK/MDPVEL28
d9FEzbRszip0Hh440+2lUXHRvOHBqLngRmjc7iFufuDtddg+Dfmsg1Dk5WYwg7j0
VDf1xCSaUe7xzu/YqCH38dtwUAylQHIIfw07e7OlcaapKh2Q2yA2CGnHIszQ6q6G
Bqym72FdjsW0VmNbA1jPzv+k1kUgzDzsvT1dR3lyTZSD6Vti+j0Jk+sKIPKybAiu
g1Qlv6tOdox2EEYseP8t+rXyiDGA+xYCIoDx9Z8TrVIQMtSFmy0niXuXNHLTMB9q
1qedHVHuP/JCYVMweShuzGV+BA9OIUYORapVumVEK0Wzw85Qj9QCADXXHhKhqfPR
18YkBoES58CdvT+Hkbw69Dg6/8Y7FjzCakjfTyLWfvbeZBwupoa/2VuVN8sA0kBK
qwJzbFz5qBywDJ4Uci5BYAKCdn/gmo5HL46jxEW87v4jSLTq0IGAaYpeRSUL8sXz
npHd5npnfxUNexcBJJE5i+JquyNw3RTIOBxqN6L2borigaHiQjV0/0UMMB2Q6pF1
DD18MCBK3b4S6iswJJdD1K3xfz7TSZDKLNNFrhWxKNeeghuBsoagMtbFWM/s/Ux4
u7kUri94FXT89ui49F9bIDdB+88nX4JNZRUvBiPwVMYD+RnAQH+Qi75v3Vhvfahv
B8PGZazbBS1nQmiHWR0oMPIj3NQbqbiWL2F4vJiWgUJqWLIpc+2W6dOuo+a93IkW
fxtyYNTUXqMhS6+yFjSFPdSd6B4V1pP+kOPrA6pquUr7mLGbh6lXqF8IQkWBZ//1
x8wSUNNPFe67dgYAZE4m4iWkaqJRKPgsfT8R78KnSJC5M1catiHrF6PuccWrk7EY
F+YvybQat7P5I0x1e+BRN7CgRCNeHayaSqNOV9O5paD6tStxFLmVjPmFJIFRzCV4
tHm0BSb4TPg63O3cfSiqP7LMUW5u2D5RCVPKjjZIZD24Bb/zIkxKf/HpsDnAU8sz
3XmR2vUHW07ck176WrOXjZ5Pw96v1tiCbv1vys0Rgp8lTyG1kbVCOrZhvqKrmlzH
XRovR7MwCNjlsHjrEW5hRVCjjRABiBcJ1u/7Pgo97u5lIlXJ+yE73gxVn5fzd/+h
6b4+1Doka9ExpaC2WSP2BXRDZBZ/a+M9Hhz/PfuQvbYlVGNAeM8ewqtUFz+OAHLM
6efxIKmwWsGL5IN98ShYAgd9QYOL0fK4AU+OtwYHSn/6yBU4JZhmvnc1XXdgTfEf
5LXsjT5zVX6WEOMf9jU5/9ogPKgvhSK+NqM/7+FXLPAts/R623TOBa/CgCRCk1NT
6r+vpP5cmCxrg427nhIFiV9jpsTlEkkBe1McJggrrCoQD/ZW57RoYXl3CH6UmKIE
yLP4GIl4XEcw8Kc2hiBK4Gs//FK5/jAo0gYL77DY9vTSeBdNgOoIh9OuRPi1wKvo
s4s+VM4K3QDhCfrd4FcBJ0YbmA9NBNXtTzWBqzUKE7Nz7TuA23lID/yuBTGDYMS4
dyUooM5r8HsvHZo/Hy+EvQbpsh1TLjg9smBnK1foPoSZprGYcsd8yfB5EutTFN36
TTFV4bAbM8p50pdizEF9FDa8aE5fLM0uNI9FuOhCyheIacyd9tqiVUQV98I54X3D
l4WoDREU/Ykl+zSO4U28JDocRzwVbqZuO9Q+DBST6S1oj+Yt2CY5wefRHYjjg1Nq
iAJNVavRLoXOGS5LJzYZN3je0uN7EHE3UD2WmH78qmjh1jANsErl+czooV9ieG2i
MKhMur0ay6MiFvxADLI2e7xMUjn1rFdfBtGVefwKdvL0/t+AnXUxFppYwtOnvVmr
UPydvpfGUYne0jBOK1Yi5FpTYxgdJVwUaTc5QD5P1uYLuIiOoh0HUnAKpuKaaawl
xrp/7Pr0xKNUnOCg3m9V4b1UFw5umcWJAFeHchfwLofPHIj0dgz4vW6jzXdM0WS6
onwWrb/BMMPzFsO9sFDuRLmG378HC4CDVLddpobu9DvRKMM+/n6f3RRCWPSnLwAO
ZMYoVYx91ObB60IXRrIaN1zSvBlSvIlQFjbc61GkQUmPe1jWA7P30QWEjczn6s7S
y+XoCz5nfOXIaBfaVD3+2BKcVdSKOiKMcQXNV/d9GzrMoQW2pLLXxCCK3lBJ/PAJ
H1xFT8l+RHnImDCxaYTeZUXQdrcQeOsi9d6w/1RLOZF3CGJE1EiiGT0ZUh7OKnwD
n3iQk7suweCfHBw/Luk/x++zHXz3fmYbXp4TLItRk1PAZAU/LtHCbwLyPLVRE8d2
13HgC1hatheTHkCCYSWjTUmeDymOsaSbDamzVJgUk/843MxcCrO+6FdldJ7cHsPT
JqrQs560wrSqxLaGQ2rcLHfDZOKqJmF3mL9LolR7Xa1gCm6vCpLTLUl21r1rhBuv
kqkhpWV+E85JF0X21DCd288zMyHZfOXmJoho7NHWrRNoyHaOlJhkAmHn5IPfqhqa
YMk8g1s2LNKCppMr0K817N1cWqE8MoYcQlP7Uteo19jieuxhqWuraXEmnjUhpIU4
8C5AoKxW4iKfIG394kodW8Nx7iZGr+nIzfhtmg1blzCcqRGHwXGi/rxX+KJviYhH
ZER2lCN3KD2x4RUltbAXhPg1mwXK7Zu5L3FFkEdO7c8BOUU6OyTYDxGegliDG5sZ
r6HyaOYerkJ1/FbU61fC3ImX7oiwK9l00c6aMCEBUw41nLtfHAywVUR+PJs8leI6
JRzGXNvDiQ2oEEtDgTd363uFqgLJzcUcIHrFgwVaSNPbpCY4G+nyDDwhj2LRTyIy
gNQOaRR6d2QTt4GhEE/Gtaz/2PjD3xi5iteD9VduGeLOsljWsTbSr2a18DwLIzTB
HR639yX6BRuHE+reT5yrht3yu1CbQVjXHcEz6jx8AKUV3h7oP3OiDEUdA7GOicv1
s5gmWN/hjvbrfUiNeMMM7GZyxuFdVV/CQJ9yVFvZ4w70cRT1ThLaa0iHNtNqdnGU
BgJX+y+Lqcc3L81zBO9Ab71tRAeiXMIzKQUD/CgxwQ3cAk9FPTeFFM02FnhqiQN6
MgO4syAjRmQXH6X9zVpFvKvuNIwfrtC7WIfbLFzdB45htsesQWhlpWXqrXBom9sb
JLS3TeecNwUrfaLx/Bma1V58ZXYrDNjNY3sBi6eBzmWHCMWlGANftvZPCeyimiqX
qQeAzjDRe2JqQsQJzFYTwLVpcYmulN61UDVMuveDxjBHQTHXGs/n4rIdCeNsHWbJ
GFFgSLqB+HdQBK1kUZuNg5YmWQtcseeqi95Kl2Lq60O46u2lf4cI3vrrMjQ1aO9c
JMoSb6CIMNIGWJexd/FUcOZIwnV+G8DFE8DsZv0+NOyCCRCtlptow0AJ8Xf52B1M
kl4c9POrQHZt8/7ibaiNgGQCy0oLTiKIQuwAv1Yey28ARTNn+eqFe/Z232IsKfAR
qjJclMxieKvczz/fmk9VUmle+wSNh5A69SWMLaHKnCkV9q1Jw+rF9VqflXqPWneq
mjOeaYGr4VahAJZ6e7KvUMB9QvXO57PN9aKZLfmjVOhY0Bk+MdXbLPFSqGmmv1N5
gcFOanAZVNzZ3m0eWD50HREfIWXKcAC6ut1hYGR7yybv6jYepcZ6xtRgF+dWslL5
3GI5vN/6nn3LRQim9KXUEjjeS+UO2p3uh0LkNck4iH15Z4xfShIpm3+xcB9WU0Ck
1Il2CZVN+y4CoyB1oUzTGa9wOgdrPm9nGoU+at7RAEezqyVlF0vjJUEP3yyknHbB
8BT1/WU/y6KDwUgk9+Fl0oJeAE2FXKsLvkv0CxBy5nBN3/FEgFeg1UXkxceCjbdR
ThHJ0zY7dqW/fnCRJrSRmk/htEcA2bguDS4Ct3JRH2quw3J95UtAepnAJb0vmXRJ
1MXeJuB+xFX8VK5Klf4LX9wyzPx3znFUdEyP2+eo+I5+9In/xBgZbnPq1LGXGVZj
BdWj9JD+Av74bH6XMyKtlCo8yc0P2Vp5uxbCIJIjP22Lt4Fjb1FSdPaSv5BZGHU6
z1ujDYwV9sCShKZbdpvZkPHH/IJQA7yQR7yLlLrrOTe9zl/2ijcj1lcgpQggCBZE
tG2wRTz9DU04ebSbxdf03ZMIFgTeoiD5uB+cVgH6u/xh/v0BtH3rNHyOjzNU7hQA
Yzf2jTfsWQyNuHMI51THAivNHEptak7ey2FbO1Nn1MUnKEWzw723OOAQXB5igTvN
AwRR4uhTe/MkeSyTpSYMi0kNUm19nae3HIwKusEZ3z1gfvqXhDhP9j9xq9j2UK7I
Z4PJjEMgvUjRUoIO3zkAvx1eOrvi/VCTTvML/mpS90DnuOzUXG+WaueWLUGJYUWT
zKryEdX/dMdOIibcEBx3bIv2Mw7TErITACu42PwxtD36sTDqXRGLgAboMsiF4E1K
2KMgkNKIIC9NnHfmzb0gbutUYPBgPnRkJcOCJOH460T8MqaE4sCa2D8Slxnsgdu5
O48PYYouaASgnouplrVfKWiyW9XlxKfCQmIutevSmbE5UL1hOVV90APPQCp/WEjY
VmGb2PFtxVvD777lQuqezQMm5agoPaQQNKvsizVFCkRH4VpmM00SRDZNNJlm9tMH
DLr2aaLqk4VUHXoe6tW0avjSXiFNcfQfhHKmOmFuXoEpVz9YXOQAivd2BD0AvXFC
ZN+Oq8loLcbcSMZmZwwhCfvSSvKG+f9L3hNy/DfRAUHodlBzSuUVgBZYZmNX8g/j
pyeYoQ+RAB+qXEZISMv80EMnXldN2WSVodM2PYOyWr2Co45+BZW5hushEfU0jDSE
EJ7RFIMSz1lIwJ17NXIbqFo2NcPDYhDN+UD7ZBTnQexZDpitsqG+nSUjw4P9z6al
sPhzll5sTQCO7frWcUHTHKP1aPxdOw8OQ2/9vtmbK+yAT+bmBBNbmJUt7pqSWGU/
uDM6LiJL0IHEef+1Zw+jvPCjQUTtb0A/atEEFimqfnlU88ygj0EHa5nQy/ZqboSb
MUquQcVXP0N0JA+5RLDsG/Shcg2k+2DBWlbr32gF5+brPZ9QOmlh/VmJrBI9jWOc
REJd5FBLM1vQQxflg38W+0gksofn4nRlJUJEftNia8QMXcKeUVoAoBezJYnuDeYn
CmKak/0P6eYYq/ptjlgVdvCp/FQkuhpj/FFfvucuXGMjl10ODD2XnjAEhvQuIX18
odbkgmqIovsPUnilny4hXghNBep6If3JUbH+Bq/dXx+A/2FklQqr0SCCRAbtlmA3
cyaXIPlSVw9obhmWm7wOKxciF/Ye/K0QGmZp/TkZde/FkIiBX5Lvs/+wTJ27dYjO
SGPy5DnZzwYP72SBeqHAu2ZbwnogzwvA5Sh4qhIOfkb+S3JQpZ00SEKMAQowpFk9
Hon/AIAfr0pQHh5Hl499k1M96TKg8p3YIswxEzCG6nlVeNZMWu62ZBZNuvRIZraq
WPB6rJhcJklD1VeZOzSctSezT/o9YT3gehmP07O6RiJ2s82syjNzPH6tJczh8jrM
98aFFkBpbtK4XIhHWayp5gMTeeZQOVEvs2xxvBzYW19KKQ1AKlKC7qY7dgLIk9IT
rhT1Q5w2bd0+cEB4eTxxr9Ldv8HJ0WastYndrAc2nkMtCaJsYKfw7TUuENoMugdf
Cn87lI7CDxCrRa7LlJVw5BvyVlAy5G1coEjua0V0Lqu9d1ozam/xzSofthM5XDED
sMVUZFABFWA7vHEqceb4YBw5eQyq0R6HOxsp0R4QOhXCpi+FQJFSFR7Zw/ODkMW6
9cNgoWcHgz+FhRyMyEO/zk5v783bbMoYaw8RutFTMnxTDLVgB9xlWP4nHSZ343Ef
E3lnuLONWxYIprOwxk9QVRk24D5m1C7WAxMjaZeCnA0jZMdE7mOlTtE7CCDQg52X
2Hh2xLWx6X9gTmqqXrv+VAyEz7rWPy9+Q85+Q/wt0b5hztlrZQv/A/hvkmiPqS2I
j+iXifGp9hQ+2JTwUTdEyeatiqxuH+2KIlN50k1ksJCMpFcCPs02yebMDYRBpfNK
QovF3Ac9rZTGC2RjthWfYqgleCO1vH2ZVRbj+35HEokVZez0rOF3aXNxZl5o2+CH
h9EAuOH9aR2ar0mUi/etTSd3Xfh8QONJPz2ssXIsCoyvDA91eAl+XGbAnOFH0EpK
3oOtUxPpEzO5dWgWAfuWRCjENeGgucE90XX5BlAcWlT5Hb9i+DiQLmdQB9QpGhwc
jV8XbMGUoJxitTBj7i3PAsEkRkC9Yhzt4PrNrlAZXlu6sFiUiEZLmay5R8X+WkvP
8jWki11DQS2fB3QWwvR9pFaM0bpcFx4jamkeYBGse/sxIGINXgjM9BgF7bJ0xSld
d5DKZ5F5st2mR35fJyWHbZ/8LwZXm6Jr71/JzfguqUguamwwvzf0iIzShH/wxP95
h8+RUKSP5HySQVWyd+fZBZpAiqdkJyaGoVdZdw7u2AkM2+6voEWwuVjl5ZWCJ/Gq
j2YaFelp/Ijttf0agXf3R4pP24WTF6wrpDRfsUwOH00R1yb7m2D37nrJiYotRpnZ
WEv1fu9U68Jgn/k7bhQrh4yJE5RHwPwW1pnVwylESEyBJL8Z6cxULvjjxSZuQucp
BGyPZmB3ALSvX/b4p28QWn8LB7Z/S+HuGVB9CqMDp339xJWF0hNZu5Fut4gHsOHS
pSYcTNcOeA6L/OITDNlgOi0k9xKkg6o7s78X3MiLcyNE0ehF7nHbgj1CI9EMIV0d
oYDrXLxR6E/x250xt221Lq1X5vb8zZDnWqx/B9Crf7eSylMj4tCpNqu2fGILnGM0
DPF6Odxo5qgExwL/b2uyOxG66R/0X8lGkdybIchIMpaomsr8kFvTBfUpEYnfHuua
KS6Az7s3z0bIMwFuWyx+3mUi9q0ZFmvGAmvt7t2Oc/8+t0J/rzpL1N7JS6k8tuaK
dz7tgknd5CDzeqohwjQVCgS4g/n+sp8+jM+RCuMzHVmB9vUppcEoj9KuEwLQ1LIU
r0p4LzvmNzduTtEXApCXIzK9QjtijGqY3XF27/usDgFEFTFCN8vfjnmVMhIfbnx+
PYOyMSPbfO6GwcxGJ04LNg3t1V6WAPyT8EYaZc9P1viG6FqsNaml5kS2oxISBBQQ
W9q0FMPwxf0Am3UrgmAsGgyRSs/B+j4ySoHvt9CoC4ViBX0Mqu3V/gt4HOfn4lqp
wpyVUVnIqTdfQzffKiucYDmzJ7Pjd3/ZWTVTZ3inSHEXagiKRVgzYNkREbgQttfv
YIAI+wLdMsMovAloYcVDnZlKf+POcI/65cAXLujGkxZLkfI62Q/Sn7RBVFEAvEz1
vmG8FdDQlMZ2QlBeKkDm3fr0Xslj1hTCgDhkUC083VGqGCC9ZScXAfvSHGefmtsn
hR5BjnIRjpc7Tu61eApbILqVi56JeG2dBCap7sPWobsFZglJQPD3HHLZRaiHgDPj
eQ67e8IYEW07T1Ngsvy5Lh4ntVyPgvgdseU0UQYUKwq9Ce5CKoAwS4PLSnRTRwcf
B4jmr9dFi4VG60QA5T7atR6jSHunPmVJn/2IoObhotp7qlEYGSyjzkLGSExP0Thw
ZwLOZToCocUryZFRii0wRkKZ/Yk5q2pKFiYwVnitBMnFAPR/DJ28K5rsSXqwQfmM
YsLWPlJawWbnQazHfNK8YzF8cnswwiF+uJXRvR8DrbYqO1BCex5dfAGpJtmnHUhc
ta70ZYwaGNsisOW4L7ocSZqB9CFEK9sWs+dpVLLGwDJE5WGYVE09agnOhIeIMuZC
l8Xq1VAnbFgrkiglv5jm7Y2CUQkBYS6yufpMblb+7RllX1HJ5e5oyY0AWsuuKi3D
lugG2CRSUXg/kEVpmz40yBRonPtJbQsVAUpN4LblTi73JHFzpAQ6jhCOLjR+VsHY
Z7YEf/3ZBWoq4wUIS7W3fG3MhzbDsYX1ddPT3mxioFHOHxsgtK4zNuRnSJQBUazJ
yuKwWVETZrK/6Z2vzp6PV6cvOkEgMMyPc26UXAdt/nroZ5t2hBGO5fL4kM4WBHP3
e1BCYNFc9LFUKlWp4vXQ8MIA83ehy2JCYRgCtQdY/I/+OmzpQyRDnynd+S4+0l0f
rAmHmjvOG2x3PG0V6Y/vn0ueYErh03SM4Wj7OhSact2SfB+0piopVVAp4Z0qEYPm
Xv9ESdCzm/m175tNV5jwhzFocPnW4RNNvDIq1y0ev6xdf4/B5smkN0scaggzUDF4
O8daQV92lnaGE9CcaKcDNsu+Ge9QUQposgFEKrwRhZa2bLxoRHxvdo/cCVT5vlPN
oKlSDGOH8dEaLNsFGKIKmuRK4X3IrpWQ0olXJAE3Rg8nUtV8Rq9ajYDH9dvbJikk
l0kVVCz0f/3sA+lUXt6G1D3e875YnkpjiApiaJ+zDhRRLBTwHo3mfN4QEiyhkNXG
VkctIhzp8IGzW53zcUXrBvNnfFH+z3WaF0Ab/2+hI1A2pznJ9+TZM2eSt3NHXdqa
UosYOGTEcpfgKvP6Of3BPA2RxzS4XsngTxVMDNgyJro/e3slypuNYeE7RnRdYdMQ
wosy+TL1OEzMnV1cyYMlWme4G98pxdaJLmtEXn7PjjJi6hIKK7rq6sRm5JkZjwok
cQX+0eRzCRw7jxJ8m0TccBkZnJnkECd9RlTLg85xtoWwCePQ4vrisameENqoQr7E
I3bg8/F7Z5HXEtBdUqWs8yydzjEVwCiRzEPrIkIngPZr3elIhCwarEOzqO5U8GEg
h/KyZWNLz0V5lXOTlVjA/zRFU8AKzAKTBauUF/3OHAx+E8zoygGurbacRf1dCyPU
E+1mhrAVK9HIcMxiMB3OWNIPCOg+mD1gghBcAZZrMcMIYu2SpRNtCYpdvxQyUlY+
hzh5pTgtCQ0Dizik1RAQomswCCVhh4EdfTrXwvbvXhcPOw+2lDe4aTGPIABjLqao
O2sUY5Sw/kcNofnqxvBSwA2fd0JmcbE38nZR8XabQYkTGEsoMnhw3aoouka9Oohy
28K9ftIZBrUGyXUGm7E0LVf8BvzcBVzY6aEDxJfRXISOr4UfbjDuncTfhd0rLZT9
sAntQDCznxAvLNIgGmr5fCohMMgnyElhsOEuSQ1g+X8hyP3pQIvki1Ljqc/oDG8h
IDmxeQHPsRabU5MDBsTYhCS1UxxLdMWvbDbI+9E148QbbJHTfxI1fZhcc9favFvw
ivFX0I21FdAVA3RtZ9VK3Wo5k1nUNCc8zQfLWinHSRxZKZLAWeSE32L2x5IxHs5b
etHYiOH6ljhf6Hmi86spy3VtDvdfTNZU/NPv9SutpCubLuVnLWH2bWGnUYRX+acZ
MxSQosrN/K5Dk8JsAXqJ/3spSuisoyY9dpvXvbKZU/uefEzywXbvKe+cFSWUTSyK
3CJsCTn8YGnOSjzlFPYBDNEIKJ9QiLKixprKhzLzck907cdaQE7PyoSPdtg0iAqk
SGy2nggT4GUHlGRhtLPkhqtij3PNkvTIuwK4WMLcVk844+6QSZIYfZPNWB7QnC/8
+uN3qpW4CCknq0dCuiY6Ti4Zzq7fCqS5RTyKJBhTGCfgizgM9H/BISDFC9pqTR6E
akiTH7SYntx8GV9EfYUwKj12fC0inbKVofplhIahYzm1KGebvI0M81FS0kv2MYlT
JnhQMQd+uWZNjTHSRwcFS0F7T6+23rDoDpi0qayAb8adBoZaQefpYJ16Q/Mrd+An
bQMv+UwINJs83OWF1hrDgxq2GCOHdWRGh6gKA+2JPwybBJSdNGZLOXYXjx5XlzIS
eTO5obflfUk06gvIC2dF6n+3aMM6Gpo5lXtw5aPvKVWrayehoWkrBXRQQ1cQpx4a
c8liZfEnEkLroZhBu3q1kapbPy/LzgjIqYCVnQthICP6cW2oEo8hHiXKDHg+8GTH
dkreFRULwmZbA3VyLCfqtK9Xso9H6KlWkYSwPSB+Lf/rsIafMy0IyP6T2odYMlpZ
N9fv13clxnWPHIj5gw4/Iv0FVbWnDbJB2GeW25O0vjKxpQBgJJfXJLaO8w00GYte
m9aDgihw/DUutxT3BeFlnj2xY737YowxgxMBPfQTuJqqtUJbF51sH192aj8tBVtU
XWTddMQzW5p0/FkyNGiNscGztbK7E0Ro1RIGqnRHAIQEJ+PXSKCeXrodF3CqCEec
B52geNGeo9Ss20+OkDgFUi8w7XrbI7n2B6DXHlo7or3m9QlE1cagv4S4V8jhF5tk
CuX5Y0irh+6epAldPzhpF9fxwfB7P4MvehUOOJ2yefojMrPE7290SLPkpRRwRICF
72tEHFNC0A6WhvnZEtmMvv5mJRM4O6gbAwW6sDhXtN41Or0OkhSF4s5ubEEtBMHK
G4vWqSReBioDLk7LfT9oMO/SPNsbynNhpzLeGXFAYOTd+zadqhYi1vAuBt1a+z/g
CciYEmMDdODKCLp03OKIWgWDr3Rbg50C4if3459ZcoaGwmJChcsgxARUaib2+eZu
FwqC8SaICAiwtFkg2hXRSYjQoxpwaZLrHVTGHdsr3jA6njRC8gqGBM6J2kIEQ2Ok
prwkNkShIL5ZTSpgxb+5KPWnGCZnXGHlax5CqWFU/MOs1Egoa+Dz3yxSEVDFpvQU
gzuu6Npmxxb9J4dSA5JTCXQV4vuABaueP3y/dCiVH76CuyFEG4oRAm/9fZtnp5r1
a+kjHQgQtUOz0qTz4oW5AFhQJHOI49qE/Bm8dduWrGu4HFYcYS1/c1fQ3A7prnGw
QXesiBFJWqO4qmGFPVTuKqJ2V95yD2EOLwL2ZW2/0npPYZRO8L8FxWANXG+FIigq
bB/Z5PRkLnAjhWStzPIH4UFej6z/7YYZh7OiKaeIXQbdLLpUiXVqyT/bGcACcaOs
Wypm87+rKqhbjVXUhFDqk1J+MKJvwlqM2pwQbtTs5qpIphNGHku83GQMm+9vFavj
Px2Kj6iUksc7rDxetbVPeMDMqjeoCWX+vy4jMoSIsHv9I/peMu8eMwsHwNZN/3CB
ebrnPJ9D6UWkESko0cTFgvYQUgLsu1iQGwCjuBYs3BAcWR4g9MDxxlFeckHXGXee
iJS6JYxUj9XsQCCYlWEO9Cc79WmNzXCK3d5ymABAp5Tvn4GpCRMqYYu7aR/UZz/L
VID/LySkADK+BxPgn4FXCOen4aUVU/uNqS5Kw1Wd5yOcxaJ9Ii4YZh3dqbY3ZDWg
Xd4GoI0g+mzgldYtDlxmq4kEY1LAJI7vZQVke2o94quUgJZlKgSVfI+PMKOr3M5O
2xdDk0Pq5rMtCAUyUJ1y8tz+Hc0IrGF+SXMgwOjEiG0xx27rKwLWozUjzNDu3ebj
rPoIpmjW+j6kL8yDrnfqMFaNQB0iQ1IdGGFMpdDPhtaq6GAvQ1/4DF9UlvIX5g/Q
UxImLeoONCUuE7g6fH8LrA6oc1+pA5XUDB/2nFLYSW8G3J5Mp5FUdZrJ7CGya5WU
0z81EMxRKogI4Vcm7NT9uerkZ/6e6jqUCSTeGEyqIBZrPVfY1cgvRFtrf1y66KPP
Ka2W2nmY3VJ2TUyj4usrb3CxnbKbIZvwUdb4d20m4M8R2RyZ4vFfMWnUVSrW0Qxp
aDOtpJzG5SOGTmzQiJkdaGrO1JAC9nORwS9ut3CzvSqFJsh5vVHJXqwpqqPHSQhf
wXo/iT/KhzQLA8bWT0xk++HQNhlQllbXKa6gBkvlBvfLRiikqAMvCP+vJN84gMwE
ACWkHTlIHV1XmVR3VqjWNtdGdaLiywYYwXp0+gP2N37RPyBTJ2rQ4rQ38amE8bVu
/XI1OXv8ycqwRxubCCivGopSzydnQpURQfTUQyHWk7nxSfgEMR7I8/Ok30G59v0K
RT0Kq4TGaP9RhPRcuk4LB/38wgntoVgqgnuQzr/hFcKsLi6hgKnLiTaxjyvtq4Os
oToWo0/u4AbZt+QGLFqGMW/9+MYQZI/8LUjE+3AmUPM2iJxAL33YZwObLfliWtB2
x/k6I2W3URB47BZ7FzAmyWMCEZPz+rMZ1XC2WIHGgzYrXWtvs6TVw8DQC5ANLbcM
mubAfWIx2/B4DBkzbfySAxU0DKtc31wCwoO/ltCdb9+8O1YYEsMtkZf2MamCiuRc
g41MZm9v125EauY3ER3hsRI05bFPU1sz696G3ctDgVgmRY8a67R1fGj4pt23lY9F
PPYtnJMV5kjk3sEgypWi1yzE4bQz8112qp0rUfA/cymIAO1j8jylPEjKVeRe7b27
TUY6nYUec/Mc6KTJ6vBIbsYYyX4SQhySrvQEoaq4uKsVF2iblfZTWPL/4Xrh4NxB
Fq/1UIrg5Qp+BloejcZGqWrQcThjl4LkP8mRQMH0ivQuzFh/JaMyryePwGHMEg4W
byXGqHJDq6RjJc6nRSRtsl8qzqYemLwEdKh0TfizT2/yC3KjQKfPCFyh5AR6eIyO
01NqfQXdD/smThsHbgzjHpDPO56mgX7kH0e8UZvYMeyIp2yxE6z/qynTGm90e/j0
oQR5fogZ62G3FU8V27chPw1Ud3lHH0+XjFUXiYZfLrSWanWSaDLW4+qvN7xBs4dR
iNV72uLtMFnAENs7uWOPd5I0FHezpD6mwSpXWj/00QmoqJab7a/XFNh6Hzpzi9S/
Dy6rS3LmOufYePmKShWYP4YkXC/K6f6EzNew2c1Jjr3MC+gFtLGlfWisHAKJPjkn
tN3vX77lSJeb9Tw2KBlERd/9cfu4qLrIj+NuBHRp/ZXEtN5qTWvQ2P5WJEpSqhJK
6/ekVWIP5xRlRppI2jBokI+ISnwFKBYO+QBZny/VIjlnKffLOOiUG0W5z7bc7z90
ImQ9lyVa+thnjz5pwt+0Qbww+lyp0bWBHmZeFt1gnhN6Gd7D6y0VgmDv5dpCS6BJ
Xu3ldmWsyT159Eiq07aoDXb3yYVNx5eq4Goz/1SlhaAGzoCxtWMbc/VhM69o/WpR
LbhqcBfcfWInjYAhzxSxYA0P+ZVg1H8EcHRvMVRG3v7Ew0vQo0k0iRJtxTTqzT4c
xpdEmy9+tgjBkmA3XJ5gepuJn6cvMQc3d+do+I4Y/fvw5G9226F4tOicTbdlMyBX
SAxs0BC+d+q2F5XBuMAHTMllXlAwgL3Q7Af4n0YkaTdAWKBn7rF9uMwEDEQ0wAuJ
a6+vctWJ48ZKHRLG2YPh8dp0OXeVD78SK5ACpwALy5o4ftCZ32P5ajEB+cZUc4Lu
z79zqkLlhGkIGOc5AD0d2EuDku6Gi5xBnZudcsJthZNwq1L2wZvk3r0uHxOTZcmD
6zhgd95y+cajDy68o4BeVPOncNYgHv99fUOxwI4YPIg225O8hWaRcexz13f09MFl
naXVzOUeHym6dOHNQbrUjIaZ1aDI42r4VccBLVc1tZTWA4B70H9tkb/gxRwWfR9F
JbziSKhFHK/FbIn33dzx5qRr0VBaNnAU63r5qY9z/rkOTR9C/euzNSiq5vn+Zx0N
Gh2ZoSkpSRle5Tp42Dqx3bha56JWhCtmVhq9vDxVMlJ/lbfCSty8Fpx3faZt3F80
dsUUm/QscEoXvJ6Dir+6nhqHbjEcIqK1ZXGX6cb5zOoW82eH1HvEdW74GWCfWVyL
M9+ehqmWcznkpg17z3wtIkxuiq3qS1HOSvMOW5DBVk4VWWrLfhVz+20/wGciWVT3
WcoKMjKDuXIls0QrQZj4sz2aro1rU2Q4KrCWkQP+5PuSLbDYXQDAU5RO4ViH+VK7
mBRbWyVmhLpVenoa2bt6Nc+ZSDrlgGeEEUVof2/pWMbFXCRzDKzD/MJF9NG74xkK
w9Tx1ncD3vTGNh65AV8H/HKgRoOTcTlss6rQATCrgVYqdGHcDxq4OfwMQ0kkA9Ea
fuLVelq1+Ql5lEr94iyezXyjBIS+NDSTGtQsJmwRfeQZAaDolN9WVtvie0HZlV0V
UxHlCCuqdmqoFnkPPQt4VIMYs2WlKIIv/r5G0HiDUy9H6l2F6lP8/UYLpiw2uhma
JiQrnMV8ET/CiO5NKdEZ9+qSWfCHqsWoUJ+/6AHlU/oob5QmoFhxpL1ULj59aeXq
W3AoyjafsY59Bg15UHg1adUDAF9tyosRXeC7vIpII+K2u9BqaEW6IMPi2iTZ6ZD/
9Jt78inQVNqyI5QqEXy76iH/sZy4Zo84wXZQABXjMazyPe1MdVnzHduxOhswZV+M
99aW5gKqslG5eqzLNAXfDIsfNe22LpI6zGtBN+cPX1oWW1xukqD36z2hU625UrWi
d+eWuknWIZV2gcF98glSDYKJIvO77Je9/RLoKQCoZhfCpzgUYJjifl7lwvvwe4Op
BXYY2Mp5+OZF4xb1XO2F3FKJImu3+fLfNpA+LC4dWGd2zCMXmVLKrnan0T+BfSvU
5VDSrvHw8ZgyUfHdHdOkQan1Stqb1dAUoNkoDK9iYnNklvLNQoj4sU9KQWJaKUX1
uCa8ksS460uNatXa/7UfOM1eDDkODP8cQIID7jSFWeb032o8fN8HZPmWnFN+3CB8
fE8ZZeBQ0B/OvhGIARNv7N76qWqzaJtTi6JefZCmqbmgVfnNaYbL4IS6tPbIInxE
R6Z2eB5aJI/mHQNYruVdeUSKYpoFEcd+7ODbNyHWVFQzgeDLP6VKzevx2sNmRo6k
dgAO7u95iFfa7dfm64rB1crL5d7FFkAsqCToL8ieaV0WKzk/NHWEmGdOFb6qGRDv
jzpT/JUnblSxx7LTDy/+C5AofdTsA3guUrNqGUqELB7e1JmgqBdpTr+OuCnZEc6c
6GeumD6DEXRHoGKwd+d+X/Opc/XtIwHXixcsLm3rY+O465S0yPPfwFuBEDQhnHP9
4hnxpolygPymoPfcQ94fxY9isld1ClJb3aqVJzkLCm4=
`pragma protect end_protected
