-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JIAMCo+pU8yhOUTkl7QvoyGqKBcdEBzQrh8/2AoVGotVWhNijOHji+tR1iHpiqneDJQIk5lMOawk
uYwil+66iKwWU2VRqAnvmdyb4PVjHg8v2+UIVnFi6uha5aB/P8MDhatjaeTfrhlEZdxVhq3HGAU/
gIECJXWDa0EBJ/TBAKTijSZuHmnMqWKYNMGzVc4nRoLCiQhBk+t8MAxonavIHwOSG/Lm46/VeEsc
UbR5wjtZH43YzE9dQ2O3He7bZCuxZF7ofzfrKUfqpnbybuR5tN6Vwlv6CxYUVBSKWnGen8SJq7zQ
IT2siHnhJqoQPayGSxHepVoWrpPJL3ezqY030g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6688)
`protect data_block
hYUJirVOeHnP23Gx3fPK0LzPeXgu+lP6ZlMrYDLGzjMxLBs0HeWBrzYv7RX8s45hCkifzgmCKmmH
k/QXWk9jPYpXkn3yQss9uvDjLGn66huf0GyhiqkthMKsD/zUdzEM08jVZqX3zH312NSG7kN9kvQK
kTXixHmvuPFzeNwyY9P69Onw2VxV9KOapGbvH29yXv50LUIBlOgztyFtjafxr2j3k3HaZ300O2ST
e5i5wTpmIjKxjDcjmgkwfZURRiogGs9Bk0O7E/rWXPypghlKxcB0V5Dg870GH1z6rSoUjPWeNyS/
EqHFvhM1B8Zsq+mF3mNV8jVLMI2CLNK+JJ9M9H5BkF3G8cJJ3F2JtpuwSPvq1By5YSZbhYqVAdfK
LsY4lqRxZsC/k3Dz5oDDqGQxXu43zPHvsSM3tHwHxABMOnszAvE688DfmpgdkjNoUbJFCBGpjBkv
5W41GIYsDuV0GunVE0LQm9zj+b7OcVM8gc2552X0GmtyDLT/eEOSFh3jLaMa7S0g1WKORUS7PJ1O
a57SRI6A8MU6vmb0LPd/tpi/HW3LcD8PtxIgslEIUH8CUVB5ZL7L91Exb7QhDv+3V4XNX5oz+UQZ
eefwHi3uFh4a2TDqyZsxgd5GaR0t/8JZH83UuCdsE/WOpXTl095MPKSXLMYHnRNQo5ruF+z/Tcz9
A+QL4KMKctsL8d8TEzx0qlqyDIb6KGbx8ohakl2dt5gH4x2OaFApzK3GV5JdBocsLmrD0OC3Qppq
XDAS7PWgWE7Lyjwi0qBk8K34JYXdtnLcXNA6KqFGwrhh5kgOlY5CnlK2R1rwaB92+xpIS0ZWm2Ud
SrWyUH+YhqYi3i77GbcPwtm/v8drywSIdrh6oIayfz5scIBxgTHwfxIKtAUVRjrb0XtHqReQ+4hv
NFearhaB74NZl9HJJJbOM2wzw6G/U6ADUUuvlRfcnE2+VRo0xo7EETkFUiQSZE0+2jmBL6x5qwD0
bZYCy8pKjPz3jTvj8CsiuSObvsuoXp5pooKc+AXL5euEQKBKBWwRnGbCieHEEEvun8MlcTCn/bdI
x40i8cmoWfmxRmNmHpA485/i24p+nKbOoNdWjUHbt2zqoCLgcTTs1SqsuImbBybT+aQM8Qy1+lT8
hzjUuBXEJsVKAzvn76Cp+UTtg6U5ot8UxG7psjGM8XbiqSQ3Sf9h06EB64gdg/rHsPLvRWoWWdR7
Xl59l3tPkefHyMaGVfbYuJIYJpyHgm00Rh/1JMkUPNQwobQkgyuzagJRXD0zKpp5mOIZBm2eXbLj
3FcFootHbGQ0vVjGsKdTeV4woDnHQwATotxdXmo7fhImXS+wwsWeGI+H7z8CXCQJYVKhw40LNW2J
AcH1bVRgofE8XUMCcNumXz9TXv9MzfO6EFydE/qFWSb4sP0gNVkLtVckPuML25KZ3jdElz4Y5sNM
jh8zqIre1FkGvgKBeg0UdfsYwmuFC+lLPwFLi7m/Bp6ioRKYrJzHGISYX3HB/kg5vqU3TeZEuv8i
iJ7NPnQrZgkHFg2oqsMbpui6E7WOYO6+Ry49LP/W2sHNozAhsA6Je7A2gFcNJYyDOfoyY28mf1A5
5eDvKXYvjKbME+k4uw2bHCloQ9zuxEwdKh19xwC3OxRaofOwJteI5W9kyigCi7VhKHknRJl/iR/0
7Q2bcAxvudocw31hjR9PrmnhYe1qT0xDw+Q4y/RQPBKgEFKbgXetO64Hg28/cxgd0Wn50f2pl1Yf
57sjTUP4wEpmCKIdK+LxrAvj5PVC+WO+RZTZzMt0NovQiF1dzrB7NXtbSPBpOVAbtZdRYjSmWTgP
/dEptyarlaGcy3eE0iMyLqTQBYhCZMOrlL1YkTHnrr3lIAr2Q8qqexEIcGM3OjVsTerZgG5jbJeS
X8ZD0eKGEauSs1fHGN0WNFyoY45zkmkpEE5VnaqmcF3sOQ6bOXjP56gm3S742w78TfFpuuBqb2ft
DlRF0+25KUVfiLegZ30x6jV8kOnID39FB9uRDslvpkn7ZPYToyJKVf4E4z2jQRodBxMvx7G03ZQN
1heowWyLUdIKWaI6O+85iHd3SBPVoZaowGpszFo/oJPeA4oMASZv5aT2AOXaD+kgd5rQxZ6LQlB9
jgNEj8A5ENey2/QsgTmy0W2XWjDPap3WnESdlmDJsGF8x0CohPzKSY2rLOaTq5r1oSmPZSmiHNCa
rXtaiJI/fjyDnvXuEicB7mAS+GHycLdRRpI0jEnqD68X04BlNJYVhmiTOWHoiy+6+Ts4MpVKYGeo
HoIsNJ9XQ31+u8Vh/tqteNXMWoxHyfEFtEVKjap/0VeIIocqUQIpTqCgHMkrRtYbKH0mpXN3Z9MR
3Lls/OGaTB9W6qSJaiH41oKLuGJJgpV7kVGcceKS7s1R1NVQXFOUEnJGFjZyGvuE5VjIZrwqsI4L
pfzsC7gSH0OI2jZdgMDfgcABDiHq+Aa4AhhlHdYH/nPD02poWrUZ5snIMvExdXMb8cbNBx58lHvT
CR5YD81KKgTCpisH2+e/xc0aHIwCf758j4H921BnoWR3u5+PiJ15IGmH5JjBN0lefWXc4ap8lEsw
BvUPVW7Psj2HlQHZRIfI1Ry4Gmpyzdv1xTRgVitzXU3nwIEnhgTAF7trFIUZzrjCJ2NknVV/Ly4p
HvAw0WtPxiYATGHb+lLNBng/5QwPq6DieuAkVfW3RbKnEsG6Pu+Y236PuYzwh4//Kte1YbOmsoHj
b1jUl9y+0guRqkLnTG6tef5x/RgPtXQtnAM6VNFmtxfhKpM8/abFROIuhrvTEiYUWzffaVijSbDj
MNAEBjRRwxVaZTyr7JQSFw7KoVJVlQrNjW1f/nl7RJqS4rdRAJLWL+tGbzWkBAm8C3gxYSmewhLP
EZ6CecNtkS456TbD8qY9EOFxTUwcyRuhTu7YoTEKZiXOG+to4poINigV9rwV/JuUURfuGrxYjUIz
zqI9X8XsBCb4sV0ruJfOvQAwo8+ttige584ILOIWLRqa1xtRDweXS3z4zYk8emMOowfYgVgdPuZG
SzbwHh2Nxk/hUfa2P+zDfJeCGjkfkyMEWgRel2bTG9FrCzCMOL/7Tkc15vVKDoEe09Q6+2nli54t
Doru+YVtfsyVpjRi/YLO3gXN2wnJB0jTWFCX0sNZjnKQkCu6cQ+EX0xy2nrEhaNAlthiZ3HsN+wW
c9ZfgwdqhpfHv9hekd4bmrF5fZ0nQbSPQne4Tx0t/CyqTezQJ7eIhqMhiK6XJ/Ms9q7fXNvOF9DV
dOcAhzl68niikcqLysRYwrbACq+nK72m5/GUq7XDdd+5/h8xr8/tCQHnxuWS5jD7FWiyoqtFoTum
pAsL5b36BQ88pxCWjewOs4d9FMgsl0aDg/90+OZz42b5gajg9fnEpQ3KdQd1eMGvsuumkZknPUwH
PHIY7HZFgu592X9yNOUd8CuRx7n1JdiywGyTeSaNT2t94NVDR2ZSzSyqN45blLHzsVj6SVPYDO8P
KOgNX1szpgn+G3hfh+K7oM1K/OVIIG+sJZnChSIJjSP21GstXvrzbp/iAQfdTfePWjkretDeDkuD
m5Mj2FbXrJIz+1noa5pMrzsKANQ+1gaKvMavyCPbtNqIjdbIJo9BwTcmJbT1tWKnPV2BrIQhp67z
VrpIZCiJz/gYYYLQJGmzds5upcozjZV9Q+puMgvAk9HqCW310/02FivUSYRHAxOBLsTMWj1K73vp
BwE0/3aVSUMHKtUuwroSeRhMQ6umlmlqISCbAF72BV2x+Ju1cOvc0jG0C0Y0EPJXR6Gb5bcVPdn6
Vv2NkwhhIXlaxCupxT/90UzGfx2xme7WF4YxDgizC958Lrk4vINRkCC+LVi1zlv5+Sb6QkVqhdy6
SL2BYkFJY1aabOSVbY/EybBTuh59D8iJBc3yCegK8V7NUu1Lv3Cqb/591hR42efFhVawlb6GOQin
qs7iVt+OfDja1JADG7SAT6va7Nea9TYNCjq5HBshSSNZm/Po71SPRWD2qCFrb0U25m+Vs9pCMzuW
QiqJOMyYrQg/Sirw+7GkKNvjaRV/cxAbWGuL/SbXsPMrGvNpnDjLC3kESP2mW/SAYmaBH05pFGYh
ryhQOX1OOKFmC86WqVR0IOBebXuyWSci1Qsvtq/vxoQSCzVwIYO1w0RsrPjP6LZjmQ+jYIl/iV4M
0skiyGeYVbcAXVrSlnufeFqezNdEd3PpxxJgkw41xiOn2hRlvX+DcGUFDvdJvsBROELUXumc4tpY
HQYWc1kdu47rV+SyY4hzCdC3Bkpr1V46ZaStKMjDClSfc8Y6u4dw+QmOT+vCIZaJGCcuWomtGOIU
fVtGGyWPYwf+oLqcckIvPWshlM6Hz5MmVkJQJWKiHpkS/oqC//3J3M7+xEoTO1+cAiWT/fJzYhdJ
L21KQCRVSpdz4itnRqeCdJIIJgzZACuAoQpPU3a6HhjXRkL45YH84MCiTzrCArLLdhEsyFTq6oY4
vX7vzums3Zsr2MppsCRcp6EvkMCqNMCjxivJJY8TnntqvIjO3VEkwABwR2CQfhMgwW+mzA5KAHPI
NARPfmSmprU+1LQmwQ9QDfRVDPjfCXSGVuv5MT1W3Xqfic18EU3Yke+5fogDOtvCc5dshuUjojjJ
lZg3kfxe15b3gwDDKmP0DjBOPgMvkoyybUUDvIWYCNtAWkGrOLqQYjDZl7IFe1l7UoTIxvymqeGE
FMU37AHmEEfru+rvP0UwhCn5pvIGLX+/XucYjFGhfh00kw5ldBy257nM+YWfixjoe8oFnSh7OVcM
xMsFOMQoX+QANVvOWPNzXZlhYF5qBA0srty1yxEfpXgTbiBJ2pDCqoBOjNweZnaOoNELilJFVSjP
/neTtL78plawjwLLpKhyxgsq+UsT64YqPl9MALXPFymezKR4AlAVc/RIgk8943Cv94z4NT2Wqfyz
Vob/sE+SPsHRLcPA+IVnfS2YSmWhJPedaPspbg9g93cplyMRzOyF/EHu2TMNRmm+PDU11tOlBtRs
TZknx08W454MWhkvj8JBLL7q0yUk4UYtvIqaMdkXEuPNGqc+VsUaeoNvHarUYOqMTczRxci9Hq2e
Ve9hup8rPCkPp1Awz+dKGW1hIP7kjfGG3vUoraeurdT2mfMtdhOIS+MvtSffEM5Rnom4RMBEDwfX
xLqrSgDL/lnf/dNVwZv9LFFjFpW2k+y2ITYi50eyWFwPCl7vSErX4V4rR0aapRsh6bAmoNrfzLlJ
EVOouL2klLNwvQkY62WxDa61ueoy/1lblCxJ0oh743FRHOwsvpS/HdUiPKt5jcVx4kaWDDwi0R2N
xEOf83RK+nZzzY1H81+LcEHnH0Sj2a4sxNwTdnHP1gpQ56LIv3a2cmws7axx8tVmFxEeWWN+FVW+
Eexj/wFVbA5XVLlqxtpInsJEOZTE50OEso7WZG8WsZKnG8iF6hz0zyUXG80Ac3ARoVyFtu4J4i4S
/XQQ89Eqr6EDqrDX7oP4kKqIvlfl2Xhtbm7+Uy9fzSDHI+Jm4/Tcg3vuXkMcyZPrYi2bkIQGnI3c
dc3SweSZnDbIKuD5VH8HTcbvrWA2HhLZMUuk+rgklzYFSws7xOxLm3dyW7LAZpEfpD7KYZyLirhc
09dsfct0cxtQwP6l38U3hOCjEn6RY+ZBjKYN8Stb57NLTFBEPhf3Bb1e466HyyaV8F3kbbcDMtfr
Rx+3VTNdLEFJQiIOz0/3vCZhWfY3quyX0FJnSHldrLEeI26ZEsryjjwKDuQn76BNnje2ShbDLgXH
Q+SWfCTdDUn/7Kq3XVj/8yRvO2vcwUzt2as7htDzqH2DaFCwhj/fgUo+dA61vnMkqTKgVW4j+Pm/
ayT/zRYi0AeHE3VeeIFqyzfDmH3EbrTpjtBHn9p+4D38wGsSW9YCzO4yZK7SRWn/+51F6NEvVcoF
AIk236TSq/GZrlFJEvh/xtfgfB8Jc2ku3T/vfhLnhGnDClaLGVRhklW6A0s3+Y19byjfwDNm7xjl
6sfKnPZxHGiZdzkjb2jJYsRfP4O219XvPIYWs/HUKDbacuoPua0JwNIW0R/7ESYedE6YYWFVqHDa
Cb+a2Fmdwx29ypoAxGCTojdsmU9egbaHbdUuO5R/lGrZC8zgl1XgAeI65xzjTorVHhS4lvwqu5d0
NcvY5L6s386iP5g9Z/w1fsPIObuBkHK7m+nyhWfIXUqXRlm9+6scFxouA5IPDKZtWeb2bOtwM7L7
5wiXawYllas4f+Fuq6TmpnxUDxRq8teSb0zrrF/7aC62beuzNTM1osFhHEmF5NUGH7t9D+2JAgWs
ip5LR8cuzClh2OqCXMPwGfoa0858YrZh12kX2UBhbrpXjmQEfbgMoL9h0TLZKPQSuazx9mOMZ8KE
8Orf/v1stI1pDSrMOH35gydXr0BwuSAostO3AE85bd3j8kp+cZZ1FP16hfux2odgGZW30WwAKOhO
/oxOhmoLXM4UHwsjyMTjbU0VJOhDDP3ejT/2zAtfG2740RxJRTQ2yGqoxRkphBAxQr16efTIgD2d
5ykElu9YaNzrFa2JbaUg1sYJ1UXCIA4Z2ROX0ee/x/2KvY0vbm/XiZaTYw6rO+v0OvSUioOsO7Yv
uaCNuHJAdDcxWz6IY8mw7Qnmm3McARquLkAKwkBEpR6LOGSSncMHuSJ8WJJvkGpDobBU4BNW5Asu
Da5SBPTrT76cwR2vVYO3y4l0xOHTS9Xct/jaPTbVcYWnJ6MJNydHHWBIjeQ4jwgnlgb81MCy42/q
wGE8qKpCASbaWaqkrQ3FcwdvVdga4rhdssONWTaCWslcqU/nKvWo8dF8CVyd/eVIEwu3ywBrvtIJ
F67pJt/xQk7Vlr2QuRgzHixder1OsQcxqASx9xVIF13LUxJ+84lnbWSIONSChgz/wSHZJwqo9+O8
ombuxkPDiFGR19PoQU4lK4s27oO9TawOxrG9fL8qeNggf2Ut3cNPtGsyfiLBkcpKXrtfZx6oT/vs
m+LBK2yrEcTk/7OV3QjdJ9Ke5uSwMlbTdGX4vIWr0hdbQLFmA50rt4oS0bgaVRA/Ud6Li6bhLkrw
B1Yg/jX/t/f8WoWK6XopcLHWxTd5Ee6Q//6mp0jKwfl7GIA2tCzi9EccQB6w826BFHxpnapIEg2J
lRLuTKloCRxIXlTqbpYabMind1JWISpScpZkn3TeJyGhUjLFXrCTDibBRgJJTJR6/oStz7t2MVcj
Jef80P08QkKBI7msiBMnaxUiEo8ftIRKrXLJJvxVLGE89jZIs0MhhA71KUcwMsrBr9h0crOCRygN
ymefrNJlQ9MVCLh+rPtGnjdaWmvjmtxWhwEvzGdOJ4WK3KoyAi0Pb3sHDZWZzaKRP0ZDADyd2dc6
SiB/79E3WOY0+zNvAd9qllOpBPShpCEptPbzbkcRiLp0g5wHq7d4APElg9IlOnyV8RYKhQJDlZlm
J+UOjFxVt04wB+chN/9C8WhmN+r3Z/8OPgCxL5V3P0FpMALXB1mbjWw09NxYgwoxW9pyguopswlz
IzEteacLeR2uwUeoVm5gYTMOkON99MQoewZSvsohzqUicR9rCMScocTFkEKXV4M0tTaoaDtQiTHI
ndybom8RJnCAJ2UUwOLSgbw8dnOYt1LvBELND4AFI6asZMSwzOn9JOxSci+3CQOtAVUaDDseau2t
K7YponskfH+fL3fWTzNM+aT+o/CN9D0LOdTEtS8wOOmvK3H6Qc9TnQ6BOgWSqtgLNanjH2Zl+Q8n
3Y5vRKEnoBegowiJGOlvOpGbbpnq5NjaMMrBleN7POxH2RfhhajeparbYmsdYw4plcWEJ9cTPTE3
dBids0uo8+/YwlKkGZq7gqnU3jD4PgJyZyVtZHAp5oCHL4uWXgVCc90X4oEVhRkppaQvWsd5sXWS
C00TlpP9tf8IPiKnVzSEdC7/ZKkv2IBOwt6NYb1fC70P/GEGICSfj206gNef56FaKqFpAyEDs8h+
pyktSd2ejrTjR/08a9IVPSIaCUe4BEzBVqGx/AhUONRV9WmgO0NZv+xGuw7x5nU9kJ2juqwOEVHy
PGU6ZTU2ufFNcvflq6FwPqPha4bs2QyGgFUnv85O52BzncDrxF2GgM+EAR6ZhfZ8LBumP26DZsN3
etzU/PydBtJl4etmeqlPp5rgkI4wRHcBBiaYBQ7NIlqlVzW6MeSqL8VdOoqT00oqi4YurLt7HJPl
tI/9lnIELOeVe/Fl2OQklan5ljJqfZXSGXJr9t3BO26MKYe429f1PdcpzajELDrr1jc147d9GtPU
dekLfgfZqOVwqcVyeNimX2gnzZr3kjCS22nbuahYrtECi7PMr/vYt+3l5+Ult8fd4GBaGCY1LUhg
ZuEow+KKZMnug3hqYk2HE0rwPE27RIXiUga3e8I9fhtP3unoWC7e2k2nniWlysYZUNoA556zrIxH
45EnaG/XC3ZyV6/H3B6ut+PoxIra62w+noHVuKm7WQ9mruicHgloaVaXKrgfeEFADrgLHMIqzA3d
Vbdel+3EMusoAGJf9dVQZ6QhS1m88eGN6/p2O67y9n5ygKOtySCKe9x2kGeomNd5rt37VuFCP9kU
Na8iNAy1gaOQhl4Yy0LlrbHK1WzrqjWO8A55JRZfzxPEP3B55xNVJj2ToXhELimBjILiRCzKuPbR
CarssWWvzthBb3xPShOwND1ddvcb9F7EdbsZxCMLuvMr/sgvI1Q1r2B7OzME0GqE0iwvpwNwGQ9P
MSHZotN2iCY2+07tJ6Eg8VAE/ghkrla+vDN3sCV7NVkdBzBfoPyB+AOpjqSpUtZ4NCpRUDoA4DO5
WUy4Ch6sx3v6ffX50e273lsrJ7K/MFCMRcd0/3C/CncuFkK/MorcaD1wQyNSh3HNPm3uD23kJt8p
mWqb2GywUQ6OaRww9GZdpg5uZg==
`protect end_protected
