��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,G�ss>ʂ�C��S��D/��mD��J���Y(�H���U��B��Z���qw0�Kǿ�(�yvE�e���>�)���L͠^����������8�4f.�`9�j8�.��ٺ�>�q��Ju�sUE�2�<4K��1Fgݬ�YxMI|+f~�?�Ԁ�;.msO0
��*OZF��0Ǽ�|#2�tц-bٶ���8fJ`^��U�B�$��~�(� a���xKX�!�u�m�T|�"���M6��zf-�`GG�.�4��a�E����d��h[-c%�K�Ê�X��p�%�ֵ�4�ϸ.�S�I��h @
�}y��(j_K	g��K4r��{��n�,�aq�3��UO}6�Zj ��Vۋ�+�۰��	ߍ_8^X��� (�SYCCt��>��o� 	��~2��b�2Έ�k���
2Os*\l���)���on�m聏3���#�w�Yg�
�+(�� &�b}T��[���	^�㕕��<7-CG�Z�����2U١�epP�v�e�qj�~J�� �w����O$&'���Q
�PK��]k��we��e�b�(gYRw��`[K�	�0y���0ȾeR�_"�
E��R����ćG��L9�5���L�@�~����u &��mR �/G-��=#y��?�0�3poZ���X�B���\�����?����W�#��B���
2dx|��Wt�Ū�a@�OL�,ވ`�ԕRK�v��9|��/k�r�P4�J�1k�IU���OU��p
���!e��X��Ϩ࣓�̖�QS~.;�Z`&�?��b���{�������Ny_���a-%@,�E��_������q�}	�`�XZ���}�I��w��en{�Y/��	V�4�h�݈�� e��LQU[~�D�n>2CA|�$�X6�|���A��WZ5��Z�K��u��B|j"���j���
�oyz�)���Uj�3r;?�s>���tlEB�T5N�d�g�DN�������Ы��"B�
�t�w����#,rS�J�)��$��y�J���y�*g1T���f|�g�<C%�n垎cC¬^+������h�fV=�g�Ϥ�y�zM*����[���o��&�r�b��J�&Xg  ,����g�������i���%����i���a
�6�"��V��fa	-7�Ah���Ya�Y��ʟ�_��օpT%�2��%"�808X�`�=��~�wk��bHWwZ�KS/0Yp�>ܯ]Ts�2q`���O�H
������F^�����C�|闍�̦�����;��EI�F����l8 37'�B*oDx��6���r���Q5��Yo�4� w��t�蕝�����F0q���?H[YWɐA��)�,�{�=�&�G���:���^1��e
/�L���g�j0����x��*-�z ���9!�A��X\�*��6���B�L����F鈈dqkѱ�ө����宁Gh��$�y�F��5���<Z O�M��h�!���9׊߿.}X%*9�ѫ���R2O�tJ���H���8[��-UyS�[�ȣ�I|�F�r�K��,hQ�K�X�c{��i���f����oIV0F�3S�Ǽ�l�}b��dA3�Ӝ)�.���H7vؼ�Y�������N�˝����ص�\����|F�#5���U��1���R�
N�:�>��6}���^Q8o� �ȢZ�(�h�F���hNB�D�TґW��t*�?�Ǥ!p�c ��} dC�Y���ɹ�cw+E��9(��U���4�!"�	;>�V�������6*�[��x�ek�����j�f�����'�T��k :��w3�~��H���J�����$��j��࣊��.���P��~��K����͜�>ku��q�ѩP&Q��'��8~�j���[۳���O&��r�������B�V77����Ip+�뢣=�{��2��o"���*r�,��3!V��U(��79�q�e4�1���ӈc]AϠn @APy�{�i��T�Ȃ����6�;��Ql�rv --}	.��x�K���JK{��#t~	�?�k���1��� (4�5��wY�rj�b8�g\{�y�5V�O&xB�x����Wj	 �l�mﯽ32��Eby���q��U�?�ފ{��pd�!��;[�n�i���/�j/ii-����1�d
�	q�&)� USi���;�g�A;�j3>P~m^�K�H��T ���P]h���^z�W�"3^����~y��M��%	17�{��RM�	E:����T��K��YjD/�A��R��A$�*Z���aw�4{��R�";�QAӡz���f�b1^Ķ�ܘ��r���g�����"��E[3��`�08�i�26�8�mѩ�~Gl����13DAW�c�yi����<����� �#�e�!�˨�\\��N���.�ֺ��?BƸ�\'�]�/�ђWգ����Zt_�5�(RG6��rr[�T����Kq�:�d�%�����by�"�}�kmW��tG�C�V�9��ʋܘ+噯����q`�5��cZ\ߵ熷�[�>F5&;��P)�|��Jb�,[�� nV�.c�|�K%��Y�-��X-R���f7�סr��|��ٯ�L���>*�bJ�.^@���טo!8�6]�^���4d�7i��:��{��M��5��+��x�)b�Ƿ������JO�3��eo6�<��&����-��N�ƀ�0���X�]&���q��
;ρ��(�7C�6A$;��s�q&Y֠��64��ѸVӦ��CՊ��� �ɭ��~r8��G�x�9|,d2��/s�����V�Д���ޱ�Oa��U6c�������������8��	|S�A^�nTI�������.��p�����}��AT|��PY�]$�G�$ R݉M�rC=�>����11�ǎT@��Ԟb�8c�GBE��}��AކF�R�^��n�N�]�B; ?@�IWc���ݸ��6�պ�jNʓ�`��*��v@�yW+�|8�{,����e�1+�J������ח�<��K�t�~Z轏L���uI!-�J{t��DbB��Í!�#w!��(M�iD�����vcngvÏ�v�_ pPHe:G٥Hh.p1��������0�̀NT�yAr`�AP�YCS�8+�ǖ�� �K��ʮۯ��A��3�-��ۖ�V�Z�
��5w)b�J��k2��t��ߧO���:��s�ud�K.2?t|̬PJ�j��t�O�?����@��tO�v�X��'�P���ȒS�����8�6p��+��4����t�`�0T�� ����V*OB��$*��7a�glq_'�S�=�����*r�5���R��ϱ�~����Y���y\  ���'����Xs<��G�0���(�b�����G�t1�����w��-�[����=.M3�?`�H�RUÌ�r�E���*��So��w��G
��4���� Y�G�/X����o����%�9\�����5��ݢ��F�m�6E�R�8�ƱB�?��p(��-���vOO}h�86ڑ���^t�=��߫�d�>�*I����$��9Ba+jv�:P�M�m<�D��5���͹T�ڗ.�`��d	ki��nF���s�H�� ��U���ݻN�������;�V���P�"^nw����ɏK�@��g�Cq��D@E���u��Ɠ�rM��짐��jx_�i�и�A�\�y�	"�E��ǒ
�)c����F��6�Y%�\�6i�b��^������iF���z����9��rEh��x�ڍT׆���h�Ж���B\�G;��g��F�4#�����z���q�n�X�Bu�����5�56�|'A݈Š��5��-uL"!4�)_�G�ɝ��^�!LmdoVṀ���y�_�u�V���Gz��)�En_��+������.�}����+��G���L���G�ض�4yL�׋�Sy�����[Ϋb^�/�j=�%���C$����݁O�����a��h�G�o����� ��ts��+�{.0��FRȲ���4��Gc�.h΅ӭlNB��{�Rk`�`u'�	6����QGf�/��.)�E�)q�e�N���_��y�сy���K(3��q�ijm��U���U��g��PDnR��ơ:S}e�L-+��"^��3'��o5bK�f�����,?f��D��DX�֯yX��5���,�"������wڬ�fE[G�dЦhpL2��ޓ���?� �i�W�oҒ1�=꬏�A������5r\�ܲ��C��g`�.t�pr��ы�X��pj;�*��|~i8U⹵��L��ђ��k��䯗�1�ľ3k�啚�J7��Rr��K�Ky�h����}��	��+�?�G�^��J*�)��}�-_�SF�)�.Q�]F���Em-�#]:l�:��!��S�Sx�8^bӑc
��ˁ���w1 	2��/���~��m���(us������ۅ��}u��&�p���T�����6����|����Sn�/�G���/�T�VsHh��6�	��,<嫛#HN�fQC��AN���:1�A��E5 ;�iՉ��;�\H�Q��$p�cC[�:�t(O�
ۼ��]� 3
�Pʂ䰩�a¢Q;Q��1��2^)V��/�sD���_�z��'!�6��kM��@� YF�=�_0��\w}������ ��"�Y����ٙ�_]ri�	��x����m�	���!���GR��g�x�����2):�Qr��*mG�]N����KP~�Ͻ��
�JR<����weOc�d�� ��&�����J(cV8���GQ�Pe����ec./*�������(��`Dg�������S���7D:2��IN�І���Ÿ�b`\��� 
��������ȯm�}$���s�2�����;\崹�����:��.���=�ȶp�e��"����#����<���)]�ls�`��f��n�4�c5�`��3�Macc�D�|�-�N%�bí�d�^ڐ@�[}��Q�8�dhZ��}&f&��s�2(��^�����ʁCh\�-:�\��-?4�1q�>P5��?���G�����9�Zh*�7&�O�t*G�1% ��IF�nb� c�v����Fȡ`C��㉝��Yx��
'��|tk�a������d�33�Ƭ�|�6���f� <�K�R[h�P����i���&n/t���zy Ϸ*k�hC>h[x<RE����}m;ru.}�S5�b?d3x
w޻:��4��N&�^:i|"P��9�S�:����5�$bo�����d7*n�U��"����R�I��6�1��D7m���,3_	4O��}w3��x���eq�{j�` {e5��k.����UZks���~٭��.���^���Gt��HS��]�V�����
�_�Y���Ѳ�� U���xL,'xh�E�:�	U�V������I��"#U�1v��ol��jnly��X��JF�9@��+XwGO�����Ga��6����I�%�5<�AW�ģ;��n���eh�y������R��tE;㚽��	����[��r�Iee�s6��ֈ+���=�%;B�΂��}�1)P9��B������9�L