// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GwvtJcpAOwiGf+n4ewC1wcbVwnO+a8GTyS7B2K9P4FUgM/KT36GDd4L+Nptbl393iAO2gquAq5TZ
CRm2ZSqenGUHwb3z03fWYw/l+7d8FOGcqaICL/bIXSI1JtUSORe3cyMAPCFN6bzoVtPb64Hl5obK
uKBq8re/VVoSk3O0Sa2sKsl2Q/yyOiW9niyM6tF5N1ufDSlyQjrNnIMhTOJdaFxtSMmG2TSb8jOk
gdsR7F3/3Bu9P9wBn0nIpY23Q6rzhItp028to+fLThtSRcc8X87RmUjZ8oKFn+3ErV3rveVkjg1e
R4sRZmihaoBRw5i9zpASEdqsAo1ZEyeZngPsOg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9024)
sGv+wKUGDZEN7zdWitkFjpRUZrEoB3KqdKUuUuHklMJgbBrZMgZfKm7FXmi51dHOqqwWjFtJP1HZ
efQRrCYHdkQ0vo/0BO4txLDkfdafZkFetj+58O81DHYeeF+ICVQZkokGH9Jm9gIsXlayfy36lSN5
WbEjn6vuhMRCX2/XmpypKG6ACWEJDk1UkeW+vAmWTneAc2FKSYxb5psa3D1izV7bwTLexmTA5ama
YZ4InKF/GHB4KVDH+fTyZOP9YSHPmpVzKBhTTN9UWv6G5StvuF2xNhp8XVwvOYxKyh8asELWgWt2
Ql1ZuIWCDvvqKFX8ChKVtsbgwZdGlriawxq9zgG/1PrWvy/qeQwQeX7AT4zLumOtotPc1STPUk0d
RHR3X3CMAGWj/PuLN8Jqf9Pa27gbwQO9fvin6tUlonXSfrAKknwoZb8a0NjyQTkLPXbvrGCWhEXi
CYwAQF1GYH3CiRyLP5fxI0vLQZXuTrv3sxtAp6/neJRg0QmEKM+d2WOFlfPe2Gdc6vrGqeL/o01+
qjqDJBjcd/qJOdXa8wZwcLwMvwwxutwgKdXiZfniJGDCNcV3NUwbrbdoDHox8owiWZNmAXuf3zM/
rDhzXAAa0oOZXwzSl4Y4hn5U+fulfmYi3Lp9f2uNFHuM0aSolcVU10wfWQdUNvLn7hHIzUgnKn6M
i8APmTMKSTlc2kRllFcS91xTF12PfH/KEka5E/UnlN9nRkTbaxWi9DpmugeavwuYEnfEEAoc6Wcw
o91XidBohIsV3YtAW5xl1/Jcz5sHxdlb1GxQV5vl8gSA3GozyN6r1tYundruXdhOmdGnL+Oipr2I
uM0SiN3dsVF7qTkHvwlYAVWEcXT3O+jeX9POMJkMPQTK5KPijRZIRsjpxcWFkux3vxmhKmTpClVZ
yco99O6kn7l0Qnqb+JcXc4DgeTCUd38UBGY87zfnG4e5gQvk8A6op6pqyxGVIX1qhrMgug4IpAh9
n4BKQvtdrWVfvuv/hm3Uitb0f5UTcOG4xGR/F7KRA8GblDPog4rNxgJ3tp0/HjZCQJWEpZhKaST/
oSvcwiWeS+GH7a2yo6AGWhfpNxwU04QmEOMYNO6lncNO/IyyiP/w3nB/gUDfd9xSJxd6slgVQI1h
wvqmNSJ3JmQlPpxmGrJr0zU8AHBahQJVL+zXrY+eoarb18KF2raDhPjJO3XsCjjeywTe2QQ9XgAp
Wp007TLDe0IHUf8FrZPNlOdtsoh+QWUUM+YfSOQ3iQYCZrZkSeQ3Zg1mrnForDWdcZ5FpbpPvlQ3
bkt83JxabKi4lmAaOi6CKArKPUdb9JVMyRmdkPStuK415cl9dhgcuappvbOdgA8aI6cy4tEXCLEr
S7p6M7PzzGMcEikEMlvw7iMv13qlhoS8FhKxv/lY7bNqzeicbPLm1gl4rjb+sARHNsBG51lT9dJ0
AA9OVhCLUJAWoJF0e/BbHk0cHGyPonYhIKnFiBCFR2qjtF0bwf/3wdFXb6qx+sbDil/IUwRnOyzx
4ptbHCN54E3C9vjyXV0tbqze6tuvkcvzZdHG3drewdie4+N+rKFiHpF2aXb5PURR39i/E/68JmWY
cKRAD+2TDpk7wkpyEyioJJvFM2WawaQkand6Jr12VOi94KrFy8YCtfsRC3jrpYRrOEppFIAZ56+a
aHTuiDGlgudY4Jb7I5MddU+puE20ATb8VW5OuyfV+mtqkCSCJF2Ltj1lpJlNx4lCmU+YKWkYgQan
c3+0qfqphGRvOBxW6lOrcAB0VQfQT3LLt0qGz9buSjPDfEhW8hXTsSVxAlT+aww+KYuBjJW1hc2S
P0/v+6AUT/A0uqVQfymFbyL4Qx99Cvkkq/wE/nVuyRFRs8qgKldpUbPjSAQL7JDu1teAWEZpjIi6
ZfIaiwRikpFX/RisISBsEqunA3mffUQwOQghXvr2zd+VP/3HPGMgPSo0W69pselss/JY9Ayft+DD
f1xYv1GISbN0e7olYOaCnmgvJ3TUdpE8xO2wNmJq05ud5gPtF1PbIo6XddSuWuYTdYwYneUGhUtf
r3PR3cZIk+5X0qAikWGhZIGLl6TBDJvOgaJmOndrf9rxdiMHOyygqJEpcRTQ7zlLcJIQcdl3w4NW
erVRGGlmWDTA0K7RC5gxoKsHtumWApYFMdOY97VplKZGw2xx1Ew3yqCqHi0TRoo2ZWdkIRVcsgIT
JPi9ueVBVbt1vyDu8tBUm5ZWzcuHgVgkh3Anpms81pO8ftfHUC8mIBfZzdOPFReAdVXmMY6+L4fb
HjFy+8tM8Q8YImFbgD0fNkdt8cpyTWSf03mTbdp5JsS9Q9WvT03FZ3wDybRgjWRtGIOfeF7rypmo
Kg5Px6UvxWA0JLN6hZY/EnEo8sxRT47PfokcTLkA3DiYS6Qq3vdpmN72CoA5s6qUF1d1QxM6U1MN
KKNTtj7pR9IbYSwFbcpgtxJkulJfTKLWNf0/MVYJT196Z10w5Jp2DjlfoAWwvrmgR216l6MqZoyT
YsXsodVnafac2GPRJIorLcRk70EXvws8ihV+T8MNcwOLcUJR7kwnuwkMLsHIZp6z899biq9S8nL3
eMustV48KeVuGntkUweOGB/+Voqv/cJ62cRGmeyhBMNdOzAadLEBd4xnpSKDvK8Tyh9TE537V8kZ
LB8JnY58F3hw9CiSM//Y5FqVolIEwDNMP02YwJd4FCIm8C702W0bihbEI+vGxVi9jSqkbrurTWU8
Dejw2YZHMvfijgNFFwguBF7I1FIOtOhg5GqMW0+XKTPyRbQBGXcaItVWSTOv2n62xfopTCxava5j
00IFN05vYyax8xAsTFCiP743upZqIytp17IK2bS7XI69U7auZn72gm9TYYABDEuhQz5IEe6jcT5p
Xi+Z9bNZuxW4x/pBxdyeoEotExZPZZ3o7PdsKhnomDLzfLzZ0cDjJ3YjbVFzlf/bUsFr+EYYoLjs
TNqZBw+RBKW+sMTgWLlbi0QXuKlyG3EtdAMwvzi/C7lLPd95/6w6xDJoJB1UFEB/2/ux6ZBDzJag
6ZifvjPZfV5zyTb0a8Az9c6ee+8qjhZGnqYeNdbwh2eRZDGIRQLBIEjLgkspiuWDZ32bnsq2OQvD
qdecZDxVcT0tE+Evrq44g00h/14cJYWrG2dWPdLjwjaTDDvsze2tWoDy/5hLqkP87MdvVyzEKhp+
lZ+Dph7qKbs/Is0DAROWgwgZQAQVq+GtQ307XYl7Lct3aFNW+2v4Ri/dZJnhWfl+wDyv2MK9FR+w
IK6GIeNInwjiGkFZAp2YIUo69YpxyyX5KJPBy+Pj0hJ9+nbrBr0xkpOMdBKRjskIiMGvVeRObjpp
WT74OeWidOzPiqgyux8sfOTdXp6ir0LKx6IcmtrO7R/pBeXIfbZ5ESeh9cCogjKiX14NWrhTp85d
skYOGK519+FjKyT1n7iZkRnNzRp1XDra/KlJuEdQq2qrln+JAu317hlkCKf+/+7+KoFORzrzAlET
Rtop49sgN46Te9EXYSZXRDc1Bs5icMI2sUJBfLAoZM4h3QLUg3aZPNm9SpHS9YkdBDPDN7sp7ruE
co5z6/PIlDJNlSFWvlWJklpA83imW9qWbK6rmUcjag1yabFpnsgV1nQfDDAQKNsgCoSd+a/eCOo6
Cjtpg+JpGh9BbxYHVY7pmqnGxWIrRb4JZlm9y8nybwM9SM1nyW4OVxM0FWfk5JgCiP0edQqNBFbc
kkQ1tU5afQ0UXkALKq2/5mRxP4uM9HVhU+SGPN0wBFF/Qb6hSYHc1Sf4EJq42nwKdDYQZ6p/4DB8
cvEepdpY9YyYoU/ugaNNKGBgu/go9gvWYxcCo+Khf+vnw3DWJRhpwPYKjs/yCGahFeE8jw7dSOQb
HDgkNXZIkpQ7XVwmog3HiW9IGgqEeJ+ItYCH1tUZmNSvcYa1f63/RG8QdlebholeLZfCGnoO4GLE
oLqKJHIQIQwx7UwwCyhBfGrHNTI8GbVFHtd6rPfqt8IOAwWuGs3gSto2KAEHKYf/LHL92y3de5aU
l4NRkHgn1WFUTIPw+1BMyKuaODW9D/ovfpR+mutb4DI9vWgwhoGeUYWiYfK8z7iCkii1cfVxcA+L
yg2H0IH5SED9Wj3OkYjhS6JwM00xvLAf8uTG1d8BphJciLfHMcTeGgIOCGBufptxdCLHH1TkiGIv
aBArzyc7dCRcAYgHAMHXfpd2ceFbUitKtsCD29Eu0SLiwnyw4vrCTDZ4o3KjNGO4jyjyRpxTiKXp
VqclxqAS51zxsDNfcmdo6KUdarWxqYIkBtTspK+09gLMZWeDwC9zf6cjnArcDlhTpBYKQLVE+Ftm
/Iu5PorwC0ghEZfjqBa3FHgVmpCcmoxxm3yhAJyc+GWuqeHIEVcZJvJhrJUnYsesGEpfnLoPxJxN
WqQGlXuuzSfwcuKoRpleep/SHl6Rk8+ZZLi7q6iXpM7qMJ7+xKZA1GkadwDAx7OXhn2o1EQQATez
rDStF6+ZAZgK79Ss+Rof8PzPeuHBqIZFubsSQWpy2YLcylj91j36LTHfIkxtN5m8KjoH0V7WMgK+
smPVSaAM/ehT0UxkJ5tuAdjh/MU8YWFnjC/RydKVtvZTVWDig63/0y1xC0wfECXfP8y6+SUa0Ias
KDTx3U1q6eEbFbVq2YpNT74VIPvSQOTf+iZQUWNPpZGGhDZmAwRUBbqzPWYmhiqa29e3Drh180ea
w9wyyp7OsPfyFyUlGTRx4c3jWBNTlUN/S13LocoPfm2NN+e/Jql9Vk+e+EUppP0OGQb1tbLlS2Km
UMReydCVk5CL2BsvVpC63wT7SK6QM3TWXZNVlQiOoDYYMyTJzvMGH8LS5zVYVqo2I5I96YqoVtC2
7VJRtHwDSPcBNBqd5jLmaOe2nGuG+wpNp7YC+KOdZmnUMJLzZEc71TPP71sEBZpn08xdRzv2l7c1
9KshDS0LTCEvBO5ITyk8vHuzErPvlmLUyRg3SYxx8Y+amtcRPVJWzxa+trvdV0aPi6ia55/p5l5S
NWOezi9twTOlJRmnDALNsEzk2NH25i8TlGYmqzDnpV2j3eOmKMc0o4nDT7Vvijf1FOlrDkHaOvhO
haHmb39URYYTapaKKTDu9XOTwwlMrQhX69bfig9IIW1FhS1Yta1226Kfs2Kacc2j/SZhiG4OkOFm
VzBXlIRVQvdjIdkXuPwaJcTFfMQEN42WPJLvinfluj/g6KrfgN/hGLksfmYtBOlSPoDPiI7PNB/r
FPxKo+VBhcOC1xfci32nQqLAIwszNL3cMDXE0bpDB7XjbRHPTqcf/mlmT1PQJ5MAQ5NepsfzjCvW
+2QN8zD/hNEr1a+pLYfSj011eP5fPeEHamkb2jlfMJEuN7QJQ4fpkQGxK8bXuWoQbTy2X4XU/bmr
8Cbljew46KhTXXCsZa5ECxNAqb03p/mYzxsRBEfIgqc/w6gelLwCsDHSCf1mrybcu2o6YeoDmKsV
S39J5/KZJ0G2f+Z2uJkHQ+VtIh+NmFDFK1/f/hdPsGHFgSBI3+6kTkMZhsCj8W+gHkH2jgk2B4fe
d2RRGB2SL94b1jzPDkzWVTTpHRrzpRm1ZEQEhOtMVWh+4b15UNdixWjF3fj7G2sHuVqxtiidvthf
H+ds4yiWAh3gDuOcDCp319NfDINhDS+zXxFgS4XXSNYFOzvkV9i9I3smRbVGdmeSPcwqY7iH5JrS
2l7U2vtNWNsktzZhOrmYY/SLn+8+eg0Wb870YhLOnvqDvLuN+W5pXJawX3MgUnmXgQBjBr+i4E4G
vB9pZz8bc2WuEmcDkVs4sA8cuGPijS2JZXomSd4lGsrfSRxL/c5mgZGEcdtty/WqYkj4nX24Q+vr
CD2efmaYFP+JGV4dIu01Jh9zFlTIVPHbnxcLyla7KYereY9IxODekE08f5gxnZXqzk9gw8WksYeh
ir/pJlgSXZmE6JtTCJhOug+BHA4NxVysXrP3Vy1yZr+106SveUSALs+G+1HRlyTV4qyBRbL1b1ez
3iscyKq/bg1VWvXMcIFJe8ZJQPima9kIjF6xfUrp1KDJzgGQIbcIfCducFwpjsjtnSojdNZcuHIY
u3CeCyR2P15drN9spZ+F34GlYy1ryhJKAPGI79H4/K8OHtrH6eWGKmA+CK5T2/o7TChGraY4Tq6U
iC8+IYMnyZr1lgsWJMpOr+fC9LFrknjv9ktVp2wPOt4lqmreF1k6uwhlpg/gRgi1QGR7rHzOHEoz
JyTgrkeN/Id6yiKpxI3Am9AKK5E+RkSC/Hfw5zfKnrEjiE80Ic3Ya7k01qkv8JKkE2XxCmNekyIk
a/i6NpSQcZ/k8fRp6UTTqjDit2eWpiAAqzRigjVa5NZoePJTCULwGSaLGJ+ONxx/kIDzekafgQsd
eIJjlhxaTMI6HHdsFOFNWcpZfrDeNVke+5tXX0pToZcy7PN/QYVp0qTQ+s8RSETJIzcNqM5mhjcT
h5nrMMCdekUYoxnMMW5Vb9UBqPsN4mBfkztDibgqhFhFKLqjpWSxN/B5dX6yMuynXq+c63vMPNv3
u1eqBZ6EDX7NL7rSN1sZ2kA6oKLuYAy38F/pYd8vRzZwTqLaQm3bHPtLtDcO4YXzsGVo8MxsRTgw
x94r1QBlLNjKKMwo24reBs8xRRAl3aoeO/pt/B3P3Xe4QEi39bC0RMtWKin2rho67ed21vPCVQNZ
/Pu05wSZA4zZ5hkG2EHBxVEWMAxFI+cDbniwuHIVQoarV3f6JXHxySbxuT3du0jIETUCjk889lto
uI84Aof3CZ4SY3MeZZZieUwMpQ7PUSA65swKXqd6DpJdab4BWbFlxM3hfFaNb4kmRvHP1v1t5dKR
eFjgWKMsBZy4qugguqZGHy2ag7Ry9OTYU5P9saMw5K/TepyU69EW2U5mcI5IFjWZVyEVihFpvk9P
46UTBQd8HVwRLoXMkmM4RrDjiRdUPmhEnXiPnyu9bdYfs41oOG9Z0Qkx3zsc2bA9VhGrKNhpw3i/
81IXKjXNYOoEjeLaVyNlb77x7GNeZQjAgiIJ7s+isSU6EFVbLfmCsek2lIhdYRZqWGSx874T0kD3
1PfcQZh7xM71sGyTsVsordRZ1TKuoCsHvlG02vWfmoEgglB9z6beaT3TtN2dMEWRk43jHLbjznK/
IcuxdFA3otCtk8N3WO/pdnWVKqV9NSe4VL63SmZgtY0Mvlf5k1vHlOILcJkMQbBTV/IirsyamMvR
LLchAMlBTRyKGD9SzuFwfhZuxU1bxKz8eVxYLPgvz3lBhdleCMpd33ii0Mt1glZ46sJlOC2+40B8
pSYurj37CiD9GSHM0k3uiz+RCgQjS7z8xK0pfxJpJo9HvsjE90l5HT6GnvQ382uOU1M5+MqfpWYm
+wEt1KDHe3DZx3bKDmohRklPyj6rm7gLjA4BHM0UB3Ibn/JUfrvMTwIezDI4iaDQkytBpLq08ANO
sJWcGnW3BmZMFosXFA4EaeW7VVZPYNxdzCAinJe0UWMPSkeByZCHDVZJJmDItyLrVHCGv6t7Pm5A
VerUWHiYRYPaURsEqOZKpdSPOdCeg0BN5cswSLu92TCDabpq9WoRP7QG4IR9DwJIxeawv1mCRjev
tkffAUOdL6SXK+2o83SHHPJ8aoXTMxIwErZMfUpELA9BUh0HHbB9J3b4Qc0S1FeSRfSNpKN6sFI6
8uewfZO+46gGwld/Hedpav+rXynfTOJtFaocBTb8Aki2A1iwJpKve6/t/vLdPV1RMDVWk73HNalT
nS9BhwF/KxSOjEPJJj5ekUo0iWUuvSdLi71WN/jhF1kYTvmaSBkONVKJgDgHKpIWUku+1qdaVp5Z
HTFLkwyJjw1GZ/xgP7nHVjLJu3SiLsO+q8enq0dZWvdxqxYQ+6aWjREm+PxDV3xNjUDelWSyDOOh
/FHji3iRHCH7y2rER6e4FtUBaPhilB4v9GhCdV9tcDJuIZVwSbzpho8WQ3qGtNU/RR0UxLvOA0/H
OdSvJJ9xn7AIiLU3MHkgAudz6kbpCPEhPlEuLjlj/znjPCfyU75jU9aoaQyUIk3cXq4b3jiMSJ2+
ecxAS9ENpXsImU7rPqp2d5oBXrfdlKT0ZQoBMTF05S72dX6w9wCzUQRKzi8G+zjOuys8rCpOtzwo
+fmdWjqrbosSMnOopemD58MaJvFsgVkzBn7seXiNNSPMMrshI4gLHkwofoSMSOBVDHBLNz5oGqCW
ZJJKBabzTHdUTqjDHfiwy5rmEwGlUvzJsQdHAjiDMLu9J2sKhIoS/UUqlSmLFP+o3p1jmqmdrRau
XPIMFvcLv6LAU0wSRGm9EPmRYzWyYyjV0Cc7e/1TFMRywGesBKsFUTBkGzdvwoO1KuMSqTPbX1Xc
7HeTpJCPYRT/xMKHCWl01IFGSY9SmiGVKLD8g6mA6HJXA20IEgQR9zUsfOiasJSB0DqclkO9YTwi
fVat3siNo+zFFk4GVVty9l4ET6rJ+xYyswHmwqIuNteNmDKXL8d7/7mX8VZyabp51QpGo2yYE1Gq
31ObrEB0sclLdhfbXOz6/haqg1DLHSK2s+InwsclylmwQ15wMLLeIQjpHM5l/hG84D9zKAcPS+ez
CUWzWpUOaaSZ/u3s1YDnkgplnAmZcaaliH5N6E/9WIE/SLNmBQv2n+eey+/Eb+YPD3e8yXO8dn3h
vadjnQrQ9S/hBH0aSXEkAYjFYC4oJY6rKVqU1sg96KJ1g/jbR6dCjHqKStltMdwDTUlzzng3G/7J
PvcMhBO417AUtNzaSgddpNUyRdb2etlryz1gaIxq6adieRSrTsAAPnJF46H4YOp1qS/SdL5NidHv
9w+mjMGlKq/DKSnuSphunGUGaejgcMJAVFiGRtXydlz8JYIG69vl38EFT+D1fRhVl+4acEszOW+C
z0dOD1eoCHw5Ep3bdL9oqDrLhGijoqEKIeF+5PK+C1Rrf7GI5KIsoT1n3JgvnnhG3VDwVU0cnNW8
TB9lqHOFtogYepXs0mHk4C+HwZ25U1wkhXFByzfj4Fu8WpGqPMXBmdzO7/yqx9scm4vQNvUo3nYU
oCFU7YzAyT72GpLM05teAPxFGhaVc0r4rD9AOcbsGnuvYzeIc9LKkxYggRq1iNOFaECxXrVP1wmo
76cfSHqaTEhxcC2TpbTc2A7imx4R8qgDQNiQs10SilEf3wmPJiUSymsVPtMFg4CfeXbXWBZnGAqj
n+FaJrwkFmstCknABRjb3WNdFa+IIWORhTCW7WI66u8vjtUEGie0kPyOEjNo8ia30Wdd9j/zlZBi
7+JC3dXmlW8EJ8yze8IQvFtihqR5CNjVllx/PAJxCK56ecIQLL7Kd2hq8x1y/ToCvQGcYz6FEtK3
Ni0EeCw/IkG6l/UkKd7fzl2JCA85xwU/tPJOE5pAPW8AYQEWAUrzRvyqqZ9zQrn2nUSPbxz2WZ8W
TEiXaeaL5r6vPKVXqUfqzos4cDMSUGGokrHofKRcRlIyIYzxgHClAsk9Qa8hYmkRTSPuIiZwAuFN
93i+Spdm+H0cCNpP68G7DSZpeLq9l5bo3ruzCZUeOFoNCGWMWGS+WtIJclM32UX4UJL92HDVfyUY
Nxo/9xNxZew61Y+4Ia4HXRsdhzhJ7/2gd2j/LZ1bKUKqwzPkwH4YG/KjCkgTWFH0e/HdCkh4vINV
q99FmylxCEBMcfZ+xmdagdl+cNMymujLmgu7ZciOc85pcZWm9ssmdu4dQT3BH3EANKyUSEg6O0lP
8c21CaCusADU08RYsPDr+Y1/pHKTrVqXBE93zZrYjUSAQz7Dcu+wo4/SrReuyN9N3wUCzKcsMjxV
FZICOihWa/7agujtEUz2gYjovkMGEM9V2M9lyaez+LrHRMHNr+o3CKuWabDx0FD0aRzhpspkfjhG
1uWpwIBHRQz7Ru8Y4gVQy52AV8rOol+6wqd+5ez02RNdZV1XCZPgA9QM2CmaXUGJNZ84PbPwxp8k
cZzsV/E2+ENxfQ/N5H7rk4FFpcFncrOB/TZs7uUBbe9a/qvpAojbqgaX24csKOxoxVUEcT9GRmIh
5BmK+Eht317uNAzDGsJMBAzC+xIz+P5V/rhv+LJqYrpPhl8eEPpzV5bKn2KHdpp65libM3Opf5Cq
iJ/k3P8CHPVJikVFCno5SSTu3nBgAqG1I9ZnesXj6gqWT1HBxOqK4Ki9CsxUzu/AHJbsWfbDs7w9
8Rju2EVItHIA5Sc6iFvPbG05cLilElyzBgmQHbLPkDxVN7Tmhs+81oBe7DqLn6rezxvK3Of2YI2r
4+MtIbkiZFEn/yBU/iGhBfziEd6AM96XInNE3nEkEjZQe5j1MW9MOQf+9Y42sH9/StgFom3JcgfU
jp+i9Qv6V3cbowWoRumPFgafbxQtBarkit/zYXK6L4VLmlGiX4vPpG4++w6N3gMTzLvDweoe4/yl
vAR0RedmUV0x7oQJhZxhdg9Xzk00/g1WRmHNd9NgbRgqM1K4X074j1v8Ci0yf6OYEEEHwyhOyfGS
bFbbvyLDLOsuVg4gPFQXF/TA6tOkqUhD9I0IXP3cUlhaXFV2bT0ttNi2BZ4B4VhvOSBQPXBtRA30
yAPmUzGotLXEHyMRAad8jGb9pEVmwx3qk0BBC6hrX9xLQE/P2R9Fu2cJbjFbUmo7Vt14U4NIBYEM
joxaVpjfJ2JRraoBkwqhPRNMkEn30Jua5UMOHTzblORWfM3wN0TQyBWW1Au6tMwsuj4X6xyGCsLW
VhlMCgxPvmk6wPn58qhCnkDMWgeAQQNc6uVnC89bLUj1iBOB90i9VfLK9MfSxh0PpNv099nKKMEj
26KR+pTmhkIGcpiZNpK/vFneiKTlvB32hMegqNfPtx13/DNgsAfOVzeT7Gguo+zFmvpKtfAs0GuK
fgdrSkPvcMji0pW7QYwYx2qpEoGHBDNvfAAK9mpjDpzLdprah1s5k4wunnvXiFTZRkdM0mCayhWE
jeTlE6/0gAsA8WSdGELE/b+jTrNSDLiI3Ewo1ooByz4ZPNgqXzwXMQvfxNshSnNBarp0pNnhf5SZ
t/BfwQ72xQ9h+6mxxQxNTVCTYAXAfr/nA7g52NGRi+RD+fnS+DFnC4b/Pgopco1kkMxWFNnJlUSc
kkFKTn02XWbpOEcl10SJlDKhr5PMWt9IKczLHjjoBVNma3HbjVXsxQzdk680qEjndNe0c9dPzkcH
cmKH4YKDAuq5Wpy0IelYA2/JMOrJ6IXiBD9quj6BzidMHK9sOKtz9zidgzljPyDkh0YfcRc4UQxi
DTCrhG+dqpGjR7seaJCJ7Vf/X8U6JZYDbE8//l/SSHnktKx42OAQ8w551+8JigXpZJhgTbp0u3BQ
k5delRIp34LoDQ01Diyukw1nmJ13GkNTKUfxU8CtweAfwIc58qGTS7vRVrc2xHM5Ga83HJ+JdJqL
0CA994VKby1sFJDrBZCiU3G1irdTFaT7Q8zlDpdqFGYgnTp+XgvpPwAKcunzupRZqKS0bik+me81
R/3mF84M/hb0ykroYTEgOOffzmVuEEZaf+j0uDjobXNFTQ1B0/RncnCOOz/viJjAf6P0aIAQJAkE
y1a925UMm7pfjj7Za91SbhJvkQsWIc6nVj+kSkHmhbrQn15eg5ovmvpOq7bxUYsGO/Sm2XO0yC45
bAMItJkrjfb+GbAEJAyzvnrKaNZ1sHu5+m6FW6czzLJxNJEKoHPRlxk5VI0iF9eCfI3lI9OFDCLc
Qr6NmSuppCHvgvohzR/hysHAmQA/8DS88fT/8u+1/ZijNk2x0fPaHhIOor35lA1tonWfZlWYcrTP
NS1ft+MAYqhi9oiBj5AdIsYSCfqIfPP8Q3o8bwfGbLi5pJnRH3Z0ngkvHJm2SgxHWKoMMIMxguV0
C156bNZGBwOkqOFdWNk3ATB5b6+53iCSZ1LnMe0NoJiviONTOlK+IJ3IDbGUXTrmMeT6VZi7ARQf
gQR7n2lBPI41QeZId1J5fVqigMIZLhG5WwbQcbtW3w2YmfKCoaOxwPEn9Cozu2inrZ9aEDaFHYK9
Cq7WEHmZ91FhqPC0YZkzj9Xa
`pragma protect end_protected
