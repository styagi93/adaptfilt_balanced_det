// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 07:05:48 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cFRMs6hqIL5ucrYlUqNnDWK6Kh3tlkGXCfGK4JtqH/tqyawzUkhp8To31Q/2//cH
U4KPi403kgI7pwEr2fQ7Tfgz0vkQ+xxbyZ6+SW0kndNKlr1lIlybDNMhjcpbn/cc
BU5vjNNWnqOMtMMxCF/fpeYzRjOX8wtG1RtA7POq2L4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9104)
7e5IRFo7Iv7BuU6G6njaW4wx1h9OfiiiWsukog0emVFudhlTU0Ky3sVDj8GK1Wgz
liTyzRCvW712+VEr/Vk9Fqlsni8eUrUhY2yk2lcWc0FNeHATYxS4UxPRZksM1WcS
oSRR4l33RVAWNnDd2qO9AXFJ18xmdNIeen4upegMfxQqY4k1FOu7J+BvPrwXUx/l
YWM/cDa2esSJxziU5mRyKiBdAJ23pX60y1A3I779QbDSTx7DWLadQ/a8gziQSvak
03V+7m5/CT2Af+XXYACOo4aZEBhj+u/9f+ezdmc3Ei7bWP1f7tz8sjHukROq7vf/
UdX2PzJsP/Ks+8uAJAODkNqgs0eqzBM1eJD0ITXxwAmwAsC0pFgVP6UEuc1YobNt
Jj6I/ecMmFZ84EAT/bqmtztbonSHzaRu7zcbKzr7YaHOGCHI3DFsWbnEq6VQpUoc
4c5wD5vokugj+LzLQGwd0n23BXOuWAD2ULF/dv41zfCUN9duETfnRSoq0jW8BDZR
q2e9ofhVZ0n5dgqp/u5fzu8q4ZMK7hGEQw+2Dp6RoDFYINCvixXfk5VBzx01gi3a
heqamSbl6oq0SKFM1lYj+5VRKiRQrXdtvLnnWHlP5SyW0cQS5IM5xaWLDVSvgSIy
1hFW9DChk8rvlVLllHJmO+1tWDmrUqkdRuo8iL629Lj5hC0vFiTT/6nfYTBfB/jQ
vQj1oK88OR92F3h7Sm/gPoRirhytmXR6BUl7rXxB+iW8I46YEl7P8GD5Vmccwd1l
w9fBgYykVtzxLlhq4YpvGHDDYIAikTnp2UE3Z7cislJZSRXqod0I7m7ROPqRC8AJ
+BEsiNFcgWKz0cfteACfOHdRlaX5i02dCjv2mfeRAtbZH0ozkvpC3UtOMVKXkLgZ
957P1cWJNxCi8hY2xFTUNiqDa/VbTlEp3aPU2fGr+k5rdptZCw/9xtnpDBN+ktJX
zrqIezvgpqJSZoE2xxhgkWuzjWqzCBB5OoNoXwvWE9St6/NhWLOE+EJ5Wlm2HwQy
3U8UFCOH/R9hc2a3OBQyXwnO8oOfrALF97Ki4XU7wjOitsJiVquyAkDhI7T+ybnd
MeNVNP/NVYRpjHary+XTEb40elG+uNvaoUROTTCoN/DicGfyUjI7e1M5xEGClNhr
tZa3Ol/DNVHW6vihDkzBg46S3/dgWL/N11RQ5K+4o3r2mS+0KJSlQoZldo2i486u
qVGdrCxn+g2i5s0d9M33DnGC3Vsg8Zi04XVBHCEXVfsOU/aoNGpA/XeYvwJ3Bjgo
ZWm4C/HN90eBvoZpiHw6XRBpfCRPaw9U71RcOUyVZJ7RtIFXVsZVAdTkNq8VzaXH
3FaMWwmXkOYUryJnoGaUnYs+hBy94/cSkhuwNAb5VXqtM32Sak0rp21fnJmvg4SM
12w9BkQejW+cY+ptse+En66bBUha4vbw9BjtyeUii3yIbURLdBaxCpQYyw4YnFn0
mC0hgNvyFibIo0j7MHXrZuJuEHfBIIU6eRheDIM4bqzzLFRP3XGRAl1pByOIWtkH
4wYDs/IJh8+UT77InPEn2+rDpD+HS/U9ElN8afJQ7YqDhP7jWUbZsPAg+lkQeFfE
5/YFgyyAlQPg6cgDU2dCy+63HL9UXgE/rCo+Viuywt4hZJ82mmHXgv4JbsmlKGRU
2dB+EfAcfeiNst537UwFj907bZcNOfB55vKIUhqHprWxF5RSa8U8pcxiAJ/iIm7X
PcXlMUtpGqNn55z96LUSsO860Eze17IJBNFv/LQ2YnZf6zjDYUR0QQzGpdfW1sdn
rZjogNaFCsMvalAAyDqmYXykU+TCCtRZxNDeiEwTlJDQD3+J/pImwvANvvFmRmGF
/Qrv1n1ZsOhgmHTW7iisZNKzq4BJU/r/Y7tm5Qca4p84zrfx16pyOHilW+8VpMz5
mU0Ne650X8Am+2KAOHbK0jQ8IIHi3/xq7TIGMjT++bSXVDXctc7Z0WThgY8k+q+Z
Muqw2C7xvgAYOO+554RORviCsqNkPiXrkjpQ4z2DXfmLiQ6MOuQGfZzoj6JzAS61
BaZNWVI2PAOeM2qArnqvBdRHMx1fH8zIlslbfyQ9Kgyifyu9c+1qDzsIHA5G/ztU
AaIjN7cGRE+IGVwV4QQj4AMr/5dzHY+Skighi+78elMMuUpiYS3+d1SLZ5gYudYV
i2PKIBTFPpUyWlJ+Y4F666LQMkDyvOtaL2kyqv+9xs3nCv9GNWCQkAKxUkIZn/lq
BR5hErEfHXAzqh7gYQTZaE1VhoRzA6pr7gXm5uAxcQB1yVdEo+96uCyVRuxTWF44
w7wHWGVEv0YcZMHsC+Fs88GOo7tXexQeRKck2/f8RssV5Rqe2B2TFPhVKHdfDqh9
WAwPhHKbhKsAyTP7tEZpxD0BWfJ61Mf+bRkHXZFKTD5tMGDd2rL8MMm8icgN6aE1
BG7mCjd80GwneVeMy/g1QIwldQtjc8w904EkAS69oUxureafHqzXiT3CMHgX0z0I
dysa/XjAqofdsWEMr4B1y1KS7Ht7YR7Na+LekrTXIxaWnD/ay6ZjrqtyeEg1tB9b
mdBDwD4u1tuk2UYqf8/V5Jbbfv69tlij0zxSlJbJG9RknNmOJh77nB4DRO17Wqcf
u2Ho0z0qNPXD0nd+5C9L/tgE2I4b1/LPwOaPGyUd3heP7GS7+c3OUqQtFM5Ty9Nr
fhzJj2ZKT0K9lB0J7W4CHy4pQcwvWpuXgbqrF0ps3Hf4k+NfS3OmEYMe6s17/Nwl
Tah04/VWGjdhLZaBAWfSus8ieDmBwOkPjWyhn0TFnYJGoI//9p39avVF6VZMI3Be
40BZj+Wy2oWxfxNZsDGsFpE/wbMFF3gD6CyuWQQNmidz3X8PMSbXEns0xcb1yh4U
4CjXJcL6QbGoXEvdSqGubT/zlqjfVSVOS192A4sckyBBkKJQIYQWuDkE3zhtD67j
O218+v59En5cll2wcMBRZ6mxqamlM/ngKKZTUXp0Z9loCdYtmNws1wFwNIMHs5Ol
flNVFNp7VT5LqmGHBAM/LrwmOnYVPheqJ4PYYYkmmAGlajeD10SEyNyMdwDSY94M
y2DDonNtUuTTHpOnjVY74PnX3jdH8e0d19DKxligCwn7iEL0H6fux7XuzGNSXsYV
Ztm3ozdpafhf9Xb7TztHWUmnku72VTFlmuJDtoYxh7Tg/o+3wP7UA7cz8seIjKCL
d/9mkrRtYX1X8GdCARNRoXTfa/kZj9dHLy9RhFsZKEvTSLUBnnRRG7RIImfsq/+O
EY+W6T9wAhuo8wCZn4yCDzXqTmiwmO+MqNN0+K76c4LQratW97q1o2HBZQTyV7IA
Lqc9OOgRkSYAE3JWehk9ZKQ4q1jxjDGFNqP/YLK9APG8MPK0MNwpWvzfyW4ZYDHJ
apyvkXl+L6QNh5VqhPldTm+ZnNZ2a/aeQB5ePdYvR7DXXar4TVIlrotL7h+hdJig
lmgFXhvW4v1Um8GAcrK029ZHoua1eYCglsUbeyUR7YbV/5jNToUvIXFdcObiGDfQ
UPNDRwB5Pl0ke8CEMDPlf8qJ8H9MGEO/o8cfU2zKoJv63Lz40XvNjd/rOHikGl2N
k6NGG6IbWShljUwMdY2HNvknA/q6YS8T8foCuzIXp63WgRTr2WxrVSWbGbC2e7Jy
F8jAb5IYflgHyjP+p4z4VaUVySfzQVQZ9PF1tfnQlEenSEbLzS0/Q5PhHr+7wHCg
zIs+I7ZX4qNRtCl0SNgyhIW5yD8iCM3Hr2HahoM1dqVoJKRC7O3oIcc3MRMT6iZH
NaRz/QxO2zJpmRdrlXc7NOkuTrF1JdT0c0U7nTPpH7tuKAwcgJo/vi01nyUH4N/f
6NNUo1Zhe/QOyIrB2nyqOg+l+vdHh+I1UZbQAP2UwQnlrtVZVvs6ynS5sh8n4VIv
BuRmel32UraRH5uN4fxEo19HRaGL0wUYCR0wGQNOpYOUFT42xXRT0gi5S2JafJKH
2sm0MLfu994xZfahRT5wXabtA83HySklDGKUzKC9W63iQpTstPoMtGz400+fpPTt
qItmYyK4AVSYwAnmH5Gun1aK/98V0l3EKdumhbLICtvfEQlnAE325gapvULFKkj8
7s8p0o+gZhtP7i5cR4YfQZdu6aIKCKLGnt+AD+lAhU4K2kSYsozB8DeGkYyUiClh
NkXH9RLjqd1JDo2aY2n6qWqmyF+5KHYs4XMcMMJF2U3HOtZvXJxFnMuDvqrdEW93
hg/EzfByWqypAQ3F3QHSWuJVBXYmkpByY+3m1UQan3cGR1zMc0tHw2MoXMODp20Y
3lobMq0cVNW7XUoLVrkBMMiJfpTgw6AXuoJtbmTV4v3d+2Q/4WYED1ezareI7D9j
cKiMoWeCtjpepOhJ5tCGE2BY/m97CkgECYfA+Hr7dc1rkfd/WStxRH8IWIviXikv
ojupUnQjI15S1hO3bC9nORZJpz3/+ligQ21yjH4bbV6352xzNYN6aSh8s4lzfQhG
rnEjlw6SAh68fOJ8MCsJoDTfe7z9qSfzREYRSsdsFcAAcfdBSd73jMrJnPL5rdB9
pAPWSu/e25/0Y/7qV0mg5UEjrUDBtaSlBj6tPU9S151pT/NEwJCBrTY3LAVxjkaZ
YTI+Zqt7waHsMEsS03jCNLGWIaWWh3Jqp+u9SElS1aYKjzg9RDYdxr/soKNI/USi
wQUeyMz06V5kOfh1sVrC7rejzK7FzX+nX5EgtaxCwIcOCCyqlYbA5VCUP//jG/vw
TF48DE+0vk54xx/TAlycOAnMHCX7Qf37OFtNikvEG5NDSFnhUWAcPk+hiusvQA5h
lJfKjplUB93NPMOhdej+fVgffOZTD2eUTqMN9q/KU6rYVVPwtn9M5zLTMm6+xZJl
XkP8v5vlpWHD/cohs6ljLDDJA07hPmtxZZLISotEOduiqgCjAa1xpbQpCD8IH9BS
HmsH1wAHixQ6OU3xJOcyegYaS4/TC93ijy6gdZQz9dP5lPxTWzvU4MpkOkO6TxYp
iXHPzP48AV58S36WtOeE5R0YFG/S0z3Pbhn5A5AE3LZekSEeJjKD1crXU4QE8HKl
UjVW7VXtsF/dbEbZlNaDJPa6wzTUwKpLWKZyEO6MrJ6kvIO4dNgNZKDzLeSCFIRe
04w86HTgaamYSrgrpHQsIrXQlSo9vVXr5pustLpv0LIpTppQvuoQRPq6/4qPoDkP
zw7Wx36ufSA5+f8YZ9cPSDwalPOUyZs97pSkiRrVHUL11zUVFhu1eEOy32XYt745
aqivN3+Z7cm1U/Les5XYYDX6GgF8hFqfyUHk/3hF8e6u8YFQeA30coacf8T9ppb0
ByhThhXopah1Wx2DkL4jtc/iB8sqqvTlxn+q836ZliWaYrn+Ipi/HS/m9eCBBn7l
9lo4VX3imTmTBFws0rFGfWLDLyi9ZABIrT4dmXnbwO63yWhKKXDlVqRNKy8e29Tw
eNyRMF8zmOMXR+nrgVVpdwYQDHa6VQ4jOuoy+qfQeujW0jqfV6Jc6UsCP3XnpVN2
mHOaORVbMy97R7ikG58La6atj0+LO2tF3LHuj7eq10AWjJxo3/fKxvkjf8p6PP+U
k53hfrNlo0ADi2bEyGVDxAoO4htdPDTJcye5mi1+3kUoGwwkbtVoOiMWVgAlZWOQ
X3hl4V7Tk0QA8eb+IkIT3ZzJChB+NMEiSJXP/FKYIY0HdbPSx6Ge6MV9bs0/cV+b
i+IAZiJJsQS1Eawvbms7/CjHf1L4aUUDcxDs5JcsFQPkMyccwNukvNpR2DWNfBny
Zb/h0dhL9VmcuhwopPIgFgToeH0r8fOASMBPR01ucBdWe14UUkBgmoHQMQt6Tdsa
iTxtyS4sImtjuEfJNsgy6cL4KYX0pMu7Fkb2RTViZJX4cwc0HSuLz3dplZNAdfjB
EAIy4oroOM7aGOWLKjzQ/emxxCZSlFMQUEww7RP148+wVg6ToDcFoY+A5yaOAZO4
UIIBkqMzfnkxTBWN83tK+TdtQuesanE0SmOnnNTGbVQhh8SjiygM8SlPClVLQhrB
t5uXK44sGcV8Bf6TXbQiMWuJED4/iLvR0RsgVm2RS1WENAMlQ7eB3OkXeEr9A9tI
FcgMuLyOUZraMAO+e0RAvdL59H5IsgGbZaVRmZA/o6wEEEVz+FwezoQKrAgkgjhx
+rd+Ld0vumXb3UrPXB62LCAShNUgSGCj7L2MAADIqbMrK/tUKRiIE3AirO7AKdfY
ZX7FycNewS7gyF5tttYRDKhNZVYDE3E5rllahD7ppZJD9ZuKAQS6JBPOdz2w/6TU
5JRP2nFbkRdHbhqjcjjhvjBHgZjqkkQ7DYD+rLPw7VUaWTFF/ac3ANmAyovAR4PV
Tpo7dUcNk/L8qgOA3g4phoFdvHl0tXx3A8WtdYepLvN3ZHAI7MBL4Sgzaahk8yyv
KpKXzPB99WcNY24B/lATqTLjfDaFyNivIlbpf/JwRAQuqArXh7G554nrQH9pVgRt
E5+RXNMMPEo9ai1DxqYXCCekek3+uzzVQ8KlaE6oOVoliwEoh17LTOQcOBfhjw5r
8uANP0wAqpMr3GG9dMMpUmaQDX2cBBBzYp9oQs8A4YHtr6qNMDWe1shuDgocZKAH
85PEsPR6N7om6Pq5d4dxLT7++PP3J+SfXg+kVci21ujbcxWr0QyRfcC+qHUnJcx4
xRMBQR31YAlNIqhU+1AZ3juG2fagvE3LfovkSeuJSK5dwmcjseueH1xTwBHQodBI
JCjeaetUbse83vGRo3fKzG+LRofOtpjuv/LFlu4TtMVpH9p8BwTIcp91HxvyKjRm
paorRJb7LjHeyZc2OSljVVZwmu7WkH6rdlnJXwUjkYp5nq9Pl0MB1mhM1WKuB2xi
JlWq2cLXlbP38MEJsZSWM4QCet7eUqg4RHpqSgkeBwNm/nToEp68fhmQf6IGNYPB
F4mmZgiqNH3PpKgfY9eokTtq87qDmAe+bvtJs3bOR4HwQ0JLxl9wmyNjThcagEF3
Ra35choudoT69B/DBs6RbEafLS0AKzfKa1Pv3LM+Vw0QFwu+VwTbRCIt5kFxcJYz
eSHfXiJVQHfegvY1Wu6eN2/+sY1XxDq3KQ2VsZQqNE6VSktY/V/1sXVVh/9mvOTJ
vyvgCnvWv4+FokwA7mYh5/i3a/FI/5EK4xZv25e/EpKAkE1ra7LV6Hc4o6siJ2Oq
hQB+ahsobl14GwNQpavk8TepDFG+L3jZJ4lrwTuyZRojGX9MHVrWRofRSN+ZY8f/
gArKgsKAMCN3Qj64AKJWNseuguR/ZclrHYMT2wXRS2eGJ50NrnyepDUS8ws8xpl+
z04KRlpgvkQLmRMQuClYykiSIZfSKl6i+MPjAFG0bcCILkcdQoyPdKiOQu2SR3D6
6vGsVYt9y5M8XmNKgmZa5nGDT44MLPFokszQLJRqfiWP/OpiysQOLsTqnVvVCeaS
UKUiGVpbnyVifIFMfilOdmJwO1/ZAni4YLMFQShqwrxVHH6pmPhKK0qjT/cwcvtJ
RxY4l5CXvYDFfOB99VbMGUSdd8zRoi2HPIdeMY0HVSnkSNwv7LMHtFLASJ6B8+lK
3XJnD2Kuqg+B+MzDBUgWaZ9Y2vI/NdauC7wl1oMIYAwLywd5F6EGZP2OIhdfs64x
TEeXAYrE859dfuDCDlzgrrsBX/RM/MtACjoGHLhd9WV48ZaQEPdHInOB8XdCZsgA
FaifByrcy1IbXb9XZKtJSy3cymGl1khGLILMkUv8UNDPIsm//dPND8Zmcw8QUUdO
/HiJmxYqORECfpxxHg7wK0D3CuyaP7YqJyTSifbjmVGlucmEM7ZHuucZNVU86NRX
GaCPO0SQJHr7IOxJe+DzPifi3H2eKYSS85097z3y8RTEpk6X4X4/LRZrdfZbRX2v
KjwdZxdJcjzw/+EjgMYrOMxJqvbREDbwmeOkUEO1gDSORUqxBcTgrkS4mTisyqhF
lVm+9ZxX5KCrbDwLVirTNjQ1HMuA/kSIrA7X0DE2WjW8h3DBFdv44HEi3Oz+XjF0
zEFF7zyDr2AhfSbm7iHidxsvCyiUFqdnU/AJZLAnWfVhlVXRl4tiHf98SjkbcrjJ
i4j/VM7mYkzZhSihPPSWl1lrgNbaidONbO85oBZLw0A5+09P7M+FRT74v6DXOZS/
EHyQK35AfkCVVbw2HDSL9VVN9E5foB8MTDbQH4Tzfc90UxS1wg6aAex1ZatUM1G+
j9wx690/67GHuxWwxKqvamu9N4y8luIKeGzOVJGgRB8NlOT779R3tdBX0KUO7qYw
Rr78pdWFM6nZXJX45iiPpGe5xH9RjuXxQrrsxnFpLBI70dAjAKsv0Qb4kl8r+fdC
KQwuxqi/lf9sLmgiknhT8aT6BJlaPkzOfgUS5qmk7RTWpfnDyHS8ZEBBj5k+9Scr
oHTFU3ZuoRPKoY8661Zq8IdyrZ0oq1Yh+JprSSZKI5iquwdj+s+Tsfrix45o4Piv
QxRvURcm01dJWQC7YChlucixBQobATtFriJqO2K6ZJE0VHcCjOvZO8I1hLOWMsNq
d7F9GIMVjICp46k36CLUZ5m66/OfrPlrjyQUkwrmKWI5J4IClwoUHpaRvnkDtyaX
X9pH+dduW9ZFGz4qlA7xN9hgdTyM00QkN18TQc9+Zbx/4D98qh+zZ2ldFCDo5mUw
SSaP8JkR/4JF6OXU1liGO0jcsbL1kDw5WDtTGqwWDo2Wj5wwop2UCLMGh72fa7AD
/yE133BRh46GHchj8oF8ul1eGAqS3N6t3Af7CBZKPY7baEpbZqD4L+ZoiwPMRLVQ
SLkiFwmzDqZpifBvX6F0ODakTloD0FtlbReLO7HymOxF5urisG32YwM7JMf0RPz/
EufWuVOODkTr3edikhx+NNLBpaTcYrAuDj9QryaH1EJeoXEeYbT7mNLQ3+W3tKM/
hAuDlrMYUIM1aJz5lmEvNPqcHHMeypaHCKJ1nRlWogvMPMKqFQTFnH6eTjX6bf1r
HQiCdd+HWldFPyYNppBqslqe2/stAW7ySV3ZOH/ko/pJKbK+VRUjbhNPJWjhs9yR
M9BBe9o89VEhzTD7QF0MxVFxdzeNgmfuyxdpABTbahdPsv/xFgxRHInJ4n4SfPSW
Cuf14YxbePCmGZyPn8DsE+V2/eNkbexYmGlOsVrdWJdsYbGFxxUmFo4xrtIW1W9x
/3+zKFPCr4TLJvo3LdUsh+kx9Mz4DcPE1lKxohm/xOyGZ0uk32aBcrFh/yu/GfxY
u29FNd6UJTeutKIu0R7aG3+Sx8hqUS9AG4SBd/A0pYJN5B/u3Ez4dQOfcMUeU2RV
luj2cNCHbHuWteuuTF+zMg7TdN0hMTE+RurjhcxuutH2GB8Vnksv5OviaPfJ//FQ
UZCS3zGuyzWc76BDbFIV7qfl6SQp14oJ+1Vm0LX6Uz8pbnV0wozMTm/dUNkJ/cPK
+4gY5jObfxsSP8HTuTSmWlEVfSJplET1yvP4RH5iqueSNOGWKf72MCmszjFdpQkG
8S9b6a2XOxusMdbfpsfdYX0aqyLdZMjH3JVWWl6zyhVK+8r1G/X7G1CoG01h++JU
QwbLbSNR+Ot4T5oXv/lo+FHRvWVoSAOswJB9Rlfyt3FWKKDnrHGdIOVmWk/tsp9V
cK66w5+xHIqRUMyEHRnEaxgxfaKn0hmAhPQNh7c8y1vgvFMrGvJ8cbDAfDQH+tlz
ScRP4B5p6fSM6hboIW6y/mBp8LFB+uRHtjanXEHt9SWC3D5EXAQFE8SVStpZIkwO
/QKdKeff1vj0UGnThQEZkIrDB9YSSFJF5Sna7PX2+QchwovYAE+KwfIi2cgnMkmv
WlztG7P/N4vH+8AlzjA+hQ/xOeXir/KlmtSAK2rQafFGcd8ZkrjvQaleH5w7s0mX
hAY1QbK3uJIg2inNl+SEaHIoaCcIty21LCyfFH833nfhjI61GSxDSKU6/YYDhFoe
wuFPIBfcMfNcSz16EPvw/qdG0MjZ4DC6i1FIJvxSrDEEACTNgXdf7WEk2UgHNzoi
Dqpt76WewmV6C/KTIZJBIZ3l8xHMpHIzw47okYiqK6j988sZOWw76NBxWmayFhhU
StL1EY4BA8DLLLM4vzldd+dySGu3yTFAXgqog7jCtGnIB96Ch+9E2t4ba+9lVi7e
AXaS1d4jl3egwRcL5LYbw3Y9QzFg50EVsHC0qkbtFcPjknqpYqbc1QqyRaqyCC2T
WbBWe6DMTwQyE/s/iVMCcBJydzV6DWknIjmBRUUsEire/mzoXTxXVgmFoOp18YSI
obaiSyU4h5JttjHA2K07kiNUDxPJCLCuvMYWHy/hL2AWcqn8QCR7ws8TTcT3oOfg
sBDa0OgD9rBNWT53j0I2H0jO89ettJbW2Hce+RXDPA6zYC6EJdB6w+un6fwoZwGH
VRd/aSDtrYEKBT57kNgc7h82itiYMhiSVLJ9k6QjMT5qcvVQUIsxK9mi0MjyO4eV
pG9HfgWL63EuC8cLTlajLY265vo5tjMX/aP7POpNVUrOH6uzwG5WvacCLkeSF5j5
3XeTkwJoD+k3dWEiqiVR96GIXjk9pCij/SCbijfjgaWwWKfR2zoZXB1lHNLDGCRT
rIJWbHktQ6gCAJ43E+5FpWQZ6D8uubB1S1uAh5k4VYfWe3Fika4ADUd2HVvw8dnd
jnzrvzjYsJWtAZRH/LW7+U1UzoidL/0c8BIapFeQEKRaYJUXf6G3EUuk1bXJEN9I
ZSUH5vINXNct+jIDc4rHVWrYO5vlmkndL6awzIqYWOD8E88ZzvgjfIRNFnf3i1qm
YX07H2nu1FYiExRClCIlybc5mjlfUhHIKuEEgyugT7JjJ4ok8SHwTLYfNhzCMSwM
1mLkMlPhJfpjUHRTp5MadklCU/zJnZ66ccAXK6CdNqR4CdTIebeD6b8vCe+1iQ3q
qX+F/n3CYbeAPFp5PVgk5HysYBPE3ZFS2gkjM9QB7ICpK39kym4s+vf9zOPQW2fo
F0mIK08c6asEKLg/3POioQ/4wOQ/v0TmN4BKE8sKK6OgIlzTPS0V2wFdAhfvoasO
qEkF2H0o3TJUrM/t/UBDPXPPsesONlc+iw4Mpy9sUzb2HJhO//kVVkv9VjEYjFO7
pdHQXtplkF4ZdMSrBzIFA7mwazYwiX6Ugfc7ujR7sA23spW9E4VOQVV29jII+/aX
CBiB59xYRI2IKnmIHVBjVJr/O5KiKCvRjikDNEsarwQHWGUtuMNqS/oyU5CnLC1o
eibeym+lW9YWFb0YeA00vYR/OJaXpPKhP89drB3UjN4DptO3gq7gbsNj2jglC2ee
ARAXnLmIY0oeb9FVu/PMZC2pPZFc4t0tRWRAR71xSngfie31xWvxbgzCO/X5f1FF
b3z1TMVakV2nJP+2MC9Zc6lx2jp8Oe8i5EOOuDGFIHKhsCUL6of7M9Iy2dODj4dg
o5cfEhrH0Do3VEaCv06r9M4r5b4ZZuiFa0zUmCv1PbUiESMdtMhsfGLb02lKBvFi
JLwVSopZaa83jli4ZvUiEwe0YZNhWNVr3GQLn9b5eFclc3I5CRSJ4aeitNBDb19M
KK3yZhgi8nRNY5+1bkRNkQLwDR9cHEJdTOeFnz0uOmc3ZR4SavC3fVOC7wqU2sZg
JzigvGT883h/0goSySRyF7uqIeVNIrghWUlJHCXz22rHMZUcNMGYn+bknsj4wqP9
5rZGEfWY/8cHQwRCl8gjJeQ3KI8+vosxJPjzI77Wb/F6K7auwbf7oDr6NsQjztzp
VJ+hbjW3bWTnqnC4+fq9bXRjiKAedTKAqoCT4glq/OgFEBa+u7kt3ZttXCN88k9v
RHgwF9bIqhoiBvuEHEQbR4HIs+pNRfmm3JZbAiKja9eh0AVH1VJ1P4S4GbGY3RCQ
oWB2z1RLzkZg2B+wjwyadJjBFlPrVi4fSFVLLHJYWJf6jC9eKXIMa+I9qYX1udul
h4P/2YJq5HasDPMo6MKd1UYjSkDzu90fJT8TA1gzV6ThaFC1bOFoy3mn3zCaNzw3
dl070yHCR/FYbnZNTJDCXq6F/WhsI2uYaGnUHTTngr3xz23QDicIRey8hNBJWR19
MRuFNzFj1yMaA9TsQUW9v5l185lrSZ8C7c0zfucsEHyQvmOyO959MOXESQd6F9Iw
sGHQFvLJYUvv4sRhjtCp8lKUe3nc6NMaxUf7rFkazr8=
`pragma protect end_protected
