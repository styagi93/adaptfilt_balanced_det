-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
cF4ZOQfxJtZNYpBGoHjvZ6qffkYT9+D3wKzWTWGgOuVH/BHzUr0cbUQAERn2F3494LHBKStHw4Sy
6m+GQy9aNBxixfcMJ3c6J3hR+5vXsRB/YE+IHoUDvNetckjEct5VoHcSarJQ9x/gCetQ8BjBVN5j
4rN4i04izBkbvD4llKPD7rV2BKH4W3zTqsOo5pumn9bcWUJvoLVps38CbMR/0ORPqKPSTrpPUMci
zQtr0UQ4n/T2/DD2tMMDXA5/YM1ThaFSSyGivwc1th2C9i9vUE5Q8hNgwniFnHYt3cmVAWNfLOAg
10/lrGUAkUC51bVHBRBeCz4Q9j3jaN5NY3K7Lw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2656)
`protect data_block
9e9lamRrxGCWAKbcBdhshk5JVa2ygRJcA7J8uSgFr2qS0Iycg1zqHqkR5bw17nwqa+bDX/RM4KaK
3so5Do6KNunxaXRAizunniaegNeZZpdlY3BRuGbQ7YefP+4gatOSNGc7rFk0wFOt5knlvLqQ4Tsw
Ya8rFb65AZfXiRmojY+zJC5LSGbzAEeioauaEMcv0f3eHVVuXuYO5F1+BgYV8xzSxoQphN6knUEV
wgrdquNzgxr/uMhqOGPWEY9LQer0ccYnS0+kBS8zNOjgWvXVn/bS+P9+TmeNn6WUiHrxEbTROWDn
XQxbsWh8dzdOKaILyLXkXzKPtUcH2QFp49XUhIsyz8Xjcw1yH3crgRh7xIbhjDrBNmWFrtIWy4gN
SX+xPh7GL66+NohrO2TnTpyAi759n1C9RBkf/ytI8nyDTg/UICkqOHBJpVN9lH2jL3/h8ag59HTL
M6sW2tiN/s/LxsoSd3xBpZW/Zjfe/F6i9H6I82aLjfW4Hx8k7l78hxUM8xthWL8fDjrv2HZU4Rcy
/6nqyq5RC235+ZnuMFZx5fjnimcdiZYmHnzSgcevcMZ1K9IU/tz0nMNH08/vCEpxm+cZ4hL6AG/L
vqJmJ5a8yxfhmZDQrc2O79oDkj1jQrJF3r52Drf90HkA6qJxj5Sh/qkMlKbj7Q60s5Z4OH7GSr/o
wt/j8fgQIpsOmCdPHORVbKuC1uTLz1ZkF2UWguqLNlAJkisiBTUWCJ0t1XuQhp7MN+nyKDZDeyT6
k5BN+sCoIdI0z1PtviOvIXQwweaCwdTVR0d984smhydqDZ+8qLAbvlBHtf4N/xr8v6pkT6FTd1Ux
qXscF9klcifY3+guhvMoUSlhNUs67/36JI2ysnENzhms6QDlba0TNKMSiHmeFEP8DFCADTZ9A5Zd
aZAj7NxIuHIxMLJTMq3pz0fa9wxDHW7nP8C3Q8jlLC8FdLpyFIMRvR8WNG14btmyUgWsw+Q+6Yre
NnRqH1TTorEP1Ix1UR32pPW/vyYFbLW6+FxzgBlYFL3lQ06XtiHMOZ4/MWOgW3PJnqI0iROLTAAO
CUsYAxgMYKzHwLF4O5HAl2Yqo1lx6mpMQyGAhEZ5RfZzGXqMUXzR7AcmmndIAf9maz+j51O1JLs2
Rmub+e+Tk3xfIWKE1CbsrGURn4ImHmLiJZwVWbwslK0dTejGLK66424dHaoT1+XZGlEY4RD9upCt
AhwxC1dvLMa2iY0l8QhoUv5X51iRzEne8LLJKEkRxqscTWbFLdojp3VaH+UyBnCewwzy+ClBQsCQ
pyRGtr7vCwQ9HUg3N/yN1YuY/1NQrgDi4gHGuyFTNYSbVzlE+IBFukMtcOxn39AnYFqM95KMpfq/
ARKA8BwrCiiP/bd/wGH0TCg9pmTPg5GIPJ85RPcvOiMt3fvg+GpcvBU+rZAKEfI1gM0I2uv/MEKO
q3l+EASWmMUc6pI23l7cmnHXJDj06rnlk2jc4bXZk5v0a0dOFeta1yVXpUmysPwBu/V1XU7Rm2Ns
wx4OwbvaUf6HRdDyXzA8XpCzqiMRUDY/fB8huVAPgdTPxOcOBe2Ad5EAyjFB4vf2QVdNbUolbN9j
dLVj3+VNiSwDAtMcyoCwN6lDWUcJxcywqYbVZ8giSTYcRlcmQwuezVPtv6KRi1BmlTUZXTlHr7oc
DK+zKCCh+vogVDBuTsXzvbWOXX4sYve6NCiQX/OqiWab4G+fzWeFuwa3Jondk/GnAD9YMnwXQg2r
0hnuzNd5fe0xSJmtRC80IkbDkm0zxLJn7jsiof3ODcivVI1bgTOPEEXNsaIhV1Dir99Ucu2JFHjV
GD5YLN5e/CVubujWoftetCVB4qUMo7GTje80Cowc9x/dNmqbrZoIyReY5fqWuI4UzHhUlLRf8K/H
Ei0eKGEP5/0MuBgqjNsBszP2LoBT/wG9UbH/+jqlbdd0BlnRm608xYEPyM29L4+odjvd7CwdLIrv
qYI+KgnNxnh6Av3Eol8iNAUg3Pfj49UZ29YXyXip3M2bH6X1rArbx0xrWc2RFoEhR05mZW0NuMlC
Xaq7w6VBphlm5HA58eeUqThC0iVkbQoZwRvJX4xp9g1vMdali/LnXwDYFQJeKQjY3mR2ysrdnIiv
XJ/0GfIrXfy+Yy849UzSzbjYPGl8FII6KT23p9NnkkBPOyuD5OFYQRnXEq0Pu6d4bUrV8l7y2owH
9A7TQLQtb9VX3+XE7IjVaNC3eE/qDaH2Fdj+/DWzjPuwm/2ffZFk4GutS+kgUiMnsYGrItcqphfn
0+eU5QI1grn2wuC7mQMdRxUHR1p+9EFTPWAX6gL5+4bMZlVpw4KJW21+ylbV75MWc8lZ9Hemetsk
vDwn+wfw2X+rLould0p8ADK4lPgJ/k10OZ1cC80TXJkyYITlAE1BBdmE2/dYljZ+hHDn+D1wW8bA
3VPShdi2HUjJ1NHTr17aoRbVr62sh0W6L3IeYgYFsgDr6k87e4RogzzRCv4yNUyBHoBenT9md6Sr
qUqPovI96ikiAZE2BVU5B1VM3tbvZKNqKMZKLeQzSgh+WlfFW5GcIwzBlGkZ2JIK6EeBvDta/VQq
YF03QPq8yObvp8OCZQh+1vTp7j0WmM3uepQG2oDHC2Q56NqLKzL3KAIKSl5dxa4DGY2f+0XKdaOn
PFwl0SW8htjKvhFGwz/VraPfdqsv6Ze+vhIxnbxw/+d8ujGBHFHa/f9XyN9ITWaPBVWBNnbOqvAS
m1Q2n6tzDJKGJYIyD/jPR0NPjF8CKxeBt3YVRDu2LTPxXXI9avCbQ8foFemHDM0d+2qKVbANRdpD
8ekfcvEUjNSU1XGPLnOawCLtiiMJd89kx50E9Wi5j9kLtj0FPUaKqmQUm6NeNJz/cbPyV3Ti2VPf
nXjoC9RK4PWcexpKOGB3ZRXG5rCP97H4yFNMaY/8Fviu9xxgLKazFdbcIedq7LrQ1vzMxxD0goSH
9QIazB9E6fzX3Cks2fBDl9Rhz9piqzdliNR5V2Ouz6155QekLr9gWpM8k5C5uzwpmNDyXi5Q8kB1
KR5ct32NRSLJi0HguGuFQzFaid+sifHAVZElDPY44osgMvEcTsRhQ/qU+HhlSbUJTcutKhkyylHq
6epZJ1dMA1kqFO/mqONpcK8VM09F0tbBV4J4/CY5+zb34/gmzrbjt6wSMt9eJLtvAt7sEfnmJV0u
Zgh8muiWbdBIVubzE3CFOlceN1tlCUO/dJapJSENwsjG/UNHDdZPm+r8z8jS+AL5Nzpcn2oUokzQ
hC0ZddCBR8UHNAc+n0jDvVoLLz0hNHWIy/cdA9Yt4nSNN60WILV7blGk84jrr80aP8CyQ4Y1pjBl
9t+2B3RMUHfYl/NmLVIYFsVTFsLhC9vNkvRuCbymidT+/4OEIiG5vNM3GdN7G2nQ6JnwEB+cfyds
itGZrlTSWDBrHEMjSI58z6N6JODqutuFPN3JdQpMXBMIij/kR4xlp6SvsQnFEdHZBAtPzIL73IKr
wkqEKlf6qltfB8k9ehnYy0nhRG5xLZmywjA6nG26p8p13Q==
`protect end_protected
